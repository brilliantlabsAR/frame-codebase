`ifndef __JISP_VH__
`define __JISP_VH__


`define USE_LATTICE_EBR


`endif // __JISP_VH__
