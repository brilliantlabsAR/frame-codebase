/*
 * This file is a part of: https://github.com/brilliantlabsAR/frame-codebase
 *
 * Authored by: Rohit Rathnam / Silicon Witchery AB (rohit@siliconwitchery.com)
 *              Raj Nakarja / Brilliant Labs Limited (raj@brilliant.xyz)
 *
 * CERN Open Hardware Licence Version 2 - Permissive
 *
 * Copyright © 2023 Brilliant Labs Limited
 */

module image_gen #(
    parameter X_RESOLUTION = 76,
    parameter Y_RESOLUTION = 76,
    parameter H_FRONT_PORCH = 152, // 2x X_RESOLUTION
    parameter H_BACK_PORCH = 167, // ~ 2.2x X_RESOLUTION
    parameter V_FRONT_PORCH = 1,
    parameter V_BACK_PORCH = 2,
    parameter H_SYNC_PULSE_WIDTH = 44,
    parameter V_SYNC_PULSE_WIDTH = 5
) (
    input logic pixel_clock_in,
    input logic reset_n_in,

    output logic [9:0] pixel_data_out,
    output logic line_valid,
    output logic frame_valid
);

logic [31:0] x_counter;
logic [31:0] y_counter;
logic [31:0] pixel_counter;

logic [9:0] mem[5927:0];

always @(posedge pixel_clock_in) begin

    if(!reset_n_in) begin

        pixel_data_out <= 0;
        line_valid <= 0;
        frame_valid <= 0;

        x_counter <= 0;
        y_counter <= 0;
        pixel_counter <= 0;

    end 

    else begin
            
        // Increment counters
        if (x_counter <= (H_SYNC_PULSE_WIDTH + H_BACK_PORCH + X_RESOLUTION + H_FRONT_PORCH)) begin
            x_counter <= x_counter + 1;
        end

        else begin
            x_counter <= 0;

            if (y_counter <= (V_SYNC_PULSE_WIDTH + V_BACK_PORCH + Y_RESOLUTION + V_FRONT_PORCH)) begin
                y_counter <= y_counter + 1;
            end

            else begin
                y_counter <= 0;
            end 

        end

        // Output line valud
        if ((x_counter >= (H_SYNC_PULSE_WIDTH + H_BACK_PORCH)) &&
            (x_counter < (H_SYNC_PULSE_WIDTH + H_BACK_PORCH + X_RESOLUTION)) &&
            (y_counter >= (V_SYNC_PULSE_WIDTH + V_BACK_PORCH)) &&
            (y_counter < (V_SYNC_PULSE_WIDTH + V_BACK_PORCH + Y_RESOLUTION))) begin
                
            line_valid <= 1;

            pixel_counter <= pixel_counter + 1;
        end

        else begin
            line_valid <= 0;
        end

        // Output frame valid
        if (y_counter >= 0 &&
            y_counter < V_SYNC_PULSE_WIDTH) begin

            frame_valid <= 0;
            pixel_counter <= 0;

        end

        else begin
            frame_valid <= 1;
        end
        
        // Output pixel
        pixel_data_out <= mem[pixel_counter];

    end

end

initial begin

    mem[0] = 'd1020;
    mem[1] = 'd1020;
    mem[2] = 'd1020;
    mem[3] = 'd1020;
    mem[4] = 'd1020;
    mem[5] = 'd1020;
    mem[6] = 'd1020;
    mem[7] = 'd1020;
    mem[8] = 'd1020;
    mem[9] = 'd1020;
    mem[10] = 'd1020;
    mem[11] = 'd1020;
    mem[12] = 'd1020;
    mem[13] = 'd1020;
    mem[14] = 'd1020;
    mem[15] = 'd1020;
    mem[16] = 'd1020;
    mem[17] = 'd1020;
    mem[18] = 'd1020;
    mem[19] = 'd1020;
    mem[20] = 'd1020;
    mem[21] = 'd1020;
    mem[22] = 'd1020;
    mem[23] = 'd1020;
    mem[24] = 'd1020;
    mem[25] = 'd1020;
    mem[26] = 'd1020;
    mem[27] = 'd1020;
    mem[28] = 'd1020;
    mem[29] = 'd1020;
    mem[30] = 'd1020;
    mem[31] = 'd1020;
    mem[32] = 'd1020;
    mem[33] = 'd1020;
    mem[34] = 'd1020;
    mem[35] = 'd1020;
    mem[36] = 'd1020;
    mem[37] = 'd1020;
    mem[38] = 'd1020;
    mem[39] = 'd1020;
    mem[40] = 'd1020;
    mem[41] = 'd1020;
    mem[42] = 'd1020;
    mem[43] = 'd1020;
    mem[44] = 'd1020;
    mem[45] = 'd1020;
    mem[46] = 'd1020;
    mem[47] = 'd1020;
    mem[48] = 'd1020;
    mem[49] = 'd1020;
    mem[50] = 'd1020;
    mem[51] = 'd1020;
    mem[52] = 'd1020;
    mem[53] = 'd1020;
    mem[54] = 'd1020;
    mem[55] = 'd1020;
    mem[56] = 'd1020;
    mem[57] = 'd1020;
    mem[58] = 'd1020;
    mem[59] = 'd1020;
    mem[60] = 'd1020;
    mem[61] = 'd1020;
    mem[62] = 'd1020;
    mem[63] = 'd1020;
    mem[64] = 'd1020;
    mem[65] = 'd1020;
    mem[66] = 'd1020;
    mem[67] = 'd1020;
    mem[68] = 'd1020;
    mem[69] = 'd1020;
    mem[70] = 'd1020;
    mem[71] = 'd1020;
    mem[72] = 'd1020;
    mem[73] = 'd1020;
    mem[74] = 'd1020;
    mem[75] = 'd1020;
    mem[76] = 'd1020;
    mem[77] = 'd1020;
    mem[78] = 'd1020;
    mem[79] = 'd1020;
    mem[80] = 'd1020;
    mem[81] = 'd1020;
    mem[82] = 'd1020;
    mem[83] = 'd1020;
    mem[84] = 'd1020;
    mem[85] = 'd1020;
    mem[86] = 'd1020;
    mem[87] = 'd1020;
    mem[88] = 'd1020;
    mem[89] = 'd1020;
    mem[90] = 'd1020;
    mem[91] = 'd1020;
    mem[92] = 'd1020;
    mem[93] = 'd1020;
    mem[94] = 'd1020;
    mem[95] = 'd1020;
    mem[96] = 'd1020;
    mem[97] = 'd1020;
    mem[98] = 'd1020;
    mem[99] = 'd1020;
    mem[100] = 'd1020;
    mem[101] = 'd1020;
    mem[102] = 'd1020;
    mem[103] = 'd1020;
    mem[104] = 'd1020;
    mem[105] = 'd1020;
    mem[106] = 'd1020;
    mem[107] = 'd1020;
    mem[108] = 'd1020;
    mem[109] = 'd1020;
    mem[110] = 'd1020;
    mem[111] = 'd1020;
    mem[112] = 'd1020;
    mem[113] = 'd1020;
    mem[114] = 'd1020;
    mem[115] = 'd1020;
    mem[116] = 'd1020;
    mem[117] = 'd1020;
    mem[118] = 'd1020;
    mem[119] = 'd1020;
    mem[120] = 'd1020;
    mem[121] = 'd1020;
    mem[122] = 'd1020;
    mem[123] = 'd1020;
    mem[124] = 'd1020;
    mem[125] = 'd1020;
    mem[126] = 'd1020;
    mem[127] = 'd1020;
    mem[128] = 'd1020;
    mem[129] = 'd1020;
    mem[130] = 'd1020;
    mem[131] = 'd1020;
    mem[132] = 'd1020;
    mem[133] = 'd1020;
    mem[134] = 'd1020;
    mem[135] = 'd1020;
    mem[136] = 'd1020;
    mem[137] = 'd1020;
    mem[138] = 'd1020;
    mem[139] = 'd1020;
    mem[140] = 'd1020;
    mem[141] = 'd1020;
    mem[142] = 'd1020;
    mem[143] = 'd1020;
    mem[144] = 'd1020;
    mem[145] = 'd1020;
    mem[146] = 'd1020;
    mem[147] = 'd1020;
    mem[148] = 'd1020;
    mem[149] = 'd1020;
    mem[150] = 'd1020;
    mem[151] = 'd1020;
    mem[152] = 'd1020;
    mem[153] = 'd1020;
    mem[154] = 'd1020;
    mem[155] = 'd1020;
    mem[156] = 'd1020;
    mem[157] = 'd1020;
    mem[158] = 'd1020;
    mem[159] = 'd1020;
    mem[160] = 'd1020;
    mem[161] = 'd1020;
    mem[162] = 'd1020;
    mem[163] = 'd1020;
    mem[164] = 'd1020;
    mem[165] = 'd1020;
    mem[166] = 'd1020;
    mem[167] = 'd1020;
    mem[168] = 'd1020;
    mem[169] = 'd1020;
    mem[170] = 'd1020;
    mem[171] = 'd1020;
    mem[172] = 'd1020;
    mem[173] = 'd1020;
    mem[174] = 'd1020;
    mem[175] = 'd1020;
    mem[176] = 'd1020;
    mem[177] = 'd1020;
    mem[178] = 'd988;
    mem[179] = 'd1000;
    mem[180] = 'd704;
    mem[181] = 'd872;
    mem[182] = 'd492;
    mem[183] = 'd804;
    mem[184] = 'd340;
    mem[185] = 'd768;
    mem[186] = 'd240;
    mem[187] = 'd748;
    mem[188] = 'd196;
    mem[189] = 'd740;
    mem[190] = 'd196;
    mem[191] = 'd740;
    mem[192] = 'd236;
    mem[193] = 'd744;
    mem[194] = 'd336;
    mem[195] = 'd764;
    mem[196] = 'd480;
    mem[197] = 'd800;
    mem[198] = 'd692;
    mem[199] = 'd868;
    mem[200] = 'd940;
    mem[201] = 'd976;
    mem[202] = 'd1020;
    mem[203] = 'd1020;
    mem[204] = 'd1020;
    mem[205] = 'd1020;
    mem[206] = 'd1020;
    mem[207] = 'd1020;
    mem[208] = 'd1020;
    mem[209] = 'd1020;
    mem[210] = 'd1020;
    mem[211] = 'd1020;
    mem[212] = 'd1020;
    mem[213] = 'd1020;
    mem[214] = 'd1020;
    mem[215] = 'd1020;
    mem[216] = 'd1020;
    mem[217] = 'd1020;
    mem[218] = 'd1020;
    mem[219] = 'd1020;
    mem[220] = 'd1020;
    mem[221] = 'd1020;
    mem[222] = 'd1020;
    mem[223] = 'd1020;
    mem[224] = 'd1020;
    mem[225] = 'd1020;
    mem[226] = 'd1020;
    mem[227] = 'd1020;
    mem[228] = 'd1020;
    mem[229] = 'd1020;
    mem[230] = 'd1020;
    mem[231] = 'd1020;
    mem[232] = 'd1020;
    mem[233] = 'd1020;
    mem[234] = 'd1020;
    mem[235] = 'd1020;
    mem[236] = 'd1020;
    mem[237] = 'd1020;
    mem[238] = 'd1020;
    mem[239] = 'd1020;
    mem[240] = 'd1020;
    mem[241] = 'd1020;
    mem[242] = 'd1020;
    mem[243] = 'd1020;
    mem[244] = 'd1020;
    mem[245] = 'd1020;
    mem[246] = 'd1020;
    mem[247] = 'd1020;
    mem[248] = 'd1020;
    mem[249] = 'd1020;
    mem[250] = 'd1020;
    mem[251] = 'd1020;
    mem[252] = 'd1020;
    mem[253] = 'd1020;
    mem[254] = 'd1000;
    mem[255] = 'd1012;
    mem[256] = 'd872;
    mem[257] = 'd1000;
    mem[258] = 'd804;
    mem[259] = 'd1000;
    mem[260] = 'd768;
    mem[261] = 'd1000;
    mem[262] = 'd748;
    mem[263] = 'd1000;
    mem[264] = 'd740;
    mem[265] = 'd1000;
    mem[266] = 'd740;
    mem[267] = 'd1000;
    mem[268] = 'd744;
    mem[269] = 'd1000;
    mem[270] = 'd764;
    mem[271] = 'd1000;
    mem[272] = 'd800;
    mem[273] = 'd1000;
    mem[274] = 'd868;
    mem[275] = 'd996;
    mem[276] = 'd976;
    mem[277] = 'd1004;
    mem[278] = 'd1020;
    mem[279] = 'd1020;
    mem[280] = 'd1020;
    mem[281] = 'd1020;
    mem[282] = 'd1020;
    mem[283] = 'd1020;
    mem[284] = 'd1020;
    mem[285] = 'd1020;
    mem[286] = 'd1020;
    mem[287] = 'd1020;
    mem[288] = 'd1020;
    mem[289] = 'd1020;
    mem[290] = 'd1020;
    mem[291] = 'd1020;
    mem[292] = 'd1020;
    mem[293] = 'd1020;
    mem[294] = 'd1020;
    mem[295] = 'd1020;
    mem[296] = 'd1020;
    mem[297] = 'd1020;
    mem[298] = 'd1020;
    mem[299] = 'd1020;
    mem[300] = 'd1020;
    mem[301] = 'd1020;
    mem[302] = 'd1020;
    mem[303] = 'd1020;
    mem[304] = 'd1020;
    mem[305] = 'd1020;
    mem[306] = 'd1020;
    mem[307] = 'd1020;
    mem[308] = 'd1020;
    mem[309] = 'd1020;
    mem[310] = 'd1020;
    mem[311] = 'd1020;
    mem[312] = 'd1020;
    mem[313] = 'd1020;
    mem[314] = 'd1020;
    mem[315] = 'd1020;
    mem[316] = 'd1020;
    mem[317] = 'd1020;
    mem[318] = 'd1020;
    mem[319] = 'd1020;
    mem[320] = 'd1020;
    mem[321] = 'd1020;
    mem[322] = 'd1020;
    mem[323] = 'd1020;
    mem[324] = 'd1020;
    mem[325] = 'd1020;
    mem[326] = 'd808;
    mem[327] = 'd912;
    mem[328] = 'd408;
    mem[329] = 'd768;
    mem[330] = 'd100;
    mem[331] = 'd696;
    mem[332] = 'd88;
    mem[333] = 'd772;
    mem[334] = 'd96;
    mem[335] = 'd828;
    mem[336] = 'd112;
    mem[337] = 'd868;
    mem[338] = 'd180;
    mem[339] = 'd900;
    mem[340] = 'd224;
    mem[341] = 'd916;
    mem[342] = 'd232;
    mem[343] = 'd916;
    mem[344] = 'd184;
    mem[345] = 'd900;
    mem[346] = 'd120;
    mem[347] = 'd868;
    mem[348] = 'd92;
    mem[349] = 'd828;
    mem[350] = 'd88;
    mem[351] = 'd776;
    mem[352] = 'd128;
    mem[353] = 'd712;
    mem[354] = 'd372;
    mem[355] = 'd752;
    mem[356] = 'd780;
    mem[357] = 'd904;
    mem[358] = 'd1012;
    mem[359] = 'd1012;
    mem[360] = 'd1020;
    mem[361] = 'd1020;
    mem[362] = 'd1020;
    mem[363] = 'd1020;
    mem[364] = 'd1020;
    mem[365] = 'd1020;
    mem[366] = 'd1020;
    mem[367] = 'd1020;
    mem[368] = 'd1020;
    mem[369] = 'd1020;
    mem[370] = 'd1020;
    mem[371] = 'd1020;
    mem[372] = 'd1020;
    mem[373] = 'd1020;
    mem[374] = 'd1020;
    mem[375] = 'd1020;
    mem[376] = 'd1020;
    mem[377] = 'd1020;
    mem[378] = 'd1020;
    mem[379] = 'd1020;
    mem[380] = 'd1020;
    mem[381] = 'd1020;
    mem[382] = 'd1020;
    mem[383] = 'd1020;
    mem[384] = 'd1020;
    mem[385] = 'd1020;
    mem[386] = 'd1020;
    mem[387] = 'd1020;
    mem[388] = 'd1020;
    mem[389] = 'd1020;
    mem[390] = 'd1020;
    mem[391] = 'd1020;
    mem[392] = 'd1020;
    mem[393] = 'd1020;
    mem[394] = 'd1020;
    mem[395] = 'd1020;
    mem[396] = 'd1020;
    mem[397] = 'd1020;
    mem[398] = 'd1020;
    mem[399] = 'd1020;
    mem[400] = 'd1020;
    mem[401] = 'd1020;
    mem[402] = 'd912;
    mem[403] = 'd996;
    mem[404] = 'd768;
    mem[405] = 'd996;
    mem[406] = 'd696;
    mem[407] = 'd1012;
    mem[408] = 'd772;
    mem[409] = 'd1020;
    mem[410] = 'd828;
    mem[411] = 'd1020;
    mem[412] = 'd868;
    mem[413] = 'd1020;
    mem[414] = 'd900;
    mem[415] = 'd1020;
    mem[416] = 'd916;
    mem[417] = 'd1020;
    mem[418] = 'd916;
    mem[419] = 'd1020;
    mem[420] = 'd900;
    mem[421] = 'd1020;
    mem[422] = 'd868;
    mem[423] = 'd1020;
    mem[424] = 'd828;
    mem[425] = 'd1020;
    mem[426] = 'd776;
    mem[427] = 'd1020;
    mem[428] = 'd712;
    mem[429] = 'd1008;
    mem[430] = 'd752;
    mem[431] = 'd996;
    mem[432] = 'd904;
    mem[433] = 'd1000;
    mem[434] = 'd1012;
    mem[435] = 'd1016;
    mem[436] = 'd1020;
    mem[437] = 'd1020;
    mem[438] = 'd1020;
    mem[439] = 'd1020;
    mem[440] = 'd1020;
    mem[441] = 'd1020;
    mem[442] = 'd1020;
    mem[443] = 'd1020;
    mem[444] = 'd1020;
    mem[445] = 'd1020;
    mem[446] = 'd1020;
    mem[447] = 'd1020;
    mem[448] = 'd1020;
    mem[449] = 'd1020;
    mem[450] = 'd1020;
    mem[451] = 'd1020;
    mem[452] = 'd1020;
    mem[453] = 'd1020;
    mem[454] = 'd1020;
    mem[455] = 'd1020;
    mem[456] = 'd1020;
    mem[457] = 'd1020;
    mem[458] = 'd1020;
    mem[459] = 'd1020;
    mem[460] = 'd1020;
    mem[461] = 'd1020;
    mem[462] = 'd1020;
    mem[463] = 'd1020;
    mem[464] = 'd1020;
    mem[465] = 'd1020;
    mem[466] = 'd1020;
    mem[467] = 'd1020;
    mem[468] = 'd1020;
    mem[469] = 'd1020;
    mem[470] = 'd1020;
    mem[471] = 'd1020;
    mem[472] = 'd1020;
    mem[473] = 'd1020;
    mem[474] = 'd868;
    mem[475] = 'd936;
    mem[476] = 'd316;
    mem[477] = 'd724;
    mem[478] = 'd52;
    mem[479] = 'd704;
    mem[480] = 'd68;
    mem[481] = 'd792;
    mem[482] = 'd164;
    mem[483] = 'd872;
    mem[484] = 'd480;
    mem[485] = 'd952;
    mem[486] = 'd704;
    mem[487] = 'd992;
    mem[488] = 'd868;
    mem[489] = 'd1012;
    mem[490] = 'd924;
    mem[491] = 'd1016;
    mem[492] = 'd940;
    mem[493] = 'd1016;
    mem[494] = 'd940;
    mem[495] = 'd1016;
    mem[496] = 'd928;
    mem[497] = 'd1016;
    mem[498] = 'd876;
    mem[499] = 'd1012;
    mem[500] = 'd736;
    mem[501] = 'd992;
    mem[502] = 'd516;
    mem[503] = 'd956;
    mem[504] = 'd228;
    mem[505] = 'd876;
    mem[506] = 'd72;
    mem[507] = 'd792;
    mem[508] = 'd64;
    mem[509] = 'd708;
    mem[510] = 'd308;
    mem[511] = 'd724;
    mem[512] = 'd824;
    mem[513] = 'd924;
    mem[514] = 'd1020;
    mem[515] = 'd1020;
    mem[516] = 'd1020;
    mem[517] = 'd1020;
    mem[518] = 'd1020;
    mem[519] = 'd1020;
    mem[520] = 'd1020;
    mem[521] = 'd1020;
    mem[522] = 'd1020;
    mem[523] = 'd1020;
    mem[524] = 'd1020;
    mem[525] = 'd1020;
    mem[526] = 'd1020;
    mem[527] = 'd1020;
    mem[528] = 'd1020;
    mem[529] = 'd1020;
    mem[530] = 'd1020;
    mem[531] = 'd1020;
    mem[532] = 'd1020;
    mem[533] = 'd1020;
    mem[534] = 'd1020;
    mem[535] = 'd1020;
    mem[536] = 'd1020;
    mem[537] = 'd1020;
    mem[538] = 'd1020;
    mem[539] = 'd1020;
    mem[540] = 'd1020;
    mem[541] = 'd1020;
    mem[542] = 'd1020;
    mem[543] = 'd1020;
    mem[544] = 'd1020;
    mem[545] = 'd1020;
    mem[546] = 'd1020;
    mem[547] = 'd1020;
    mem[548] = 'd1020;
    mem[549] = 'd1020;
    mem[550] = 'd936;
    mem[551] = 'd996;
    mem[552] = 'd724;
    mem[553] = 'd996;
    mem[554] = 'd704;
    mem[555] = 'd1020;
    mem[556] = 'd792;
    mem[557] = 'd1020;
    mem[558] = 'd872;
    mem[559] = 'd1020;
    mem[560] = 'd952;
    mem[561] = 'd1020;
    mem[562] = 'd992;
    mem[563] = 'd1020;
    mem[564] = 'd1012;
    mem[565] = 'd1020;
    mem[566] = 'd1016;
    mem[567] = 'd1020;
    mem[568] = 'd1016;
    mem[569] = 'd1020;
    mem[570] = 'd1016;
    mem[571] = 'd1020;
    mem[572] = 'd1016;
    mem[573] = 'd1020;
    mem[574] = 'd1012;
    mem[575] = 'd1020;
    mem[576] = 'd992;
    mem[577] = 'd1020;
    mem[578] = 'd956;
    mem[579] = 'd1020;
    mem[580] = 'd876;
    mem[581] = 'd1020;
    mem[582] = 'd792;
    mem[583] = 'd1020;
    mem[584] = 'd708;
    mem[585] = 'd1016;
    mem[586] = 'd724;
    mem[587] = 'd996;
    mem[588] = 'd924;
    mem[589] = 'd1000;
    mem[590] = 'd1020;
    mem[591] = 'd1020;
    mem[592] = 'd1020;
    mem[593] = 'd1020;
    mem[594] = 'd1020;
    mem[595] = 'd1020;
    mem[596] = 'd1020;
    mem[597] = 'd1020;
    mem[598] = 'd1020;
    mem[599] = 'd1020;
    mem[600] = 'd1020;
    mem[601] = 'd1020;
    mem[602] = 'd1020;
    mem[603] = 'd1020;
    mem[604] = 'd1020;
    mem[605] = 'd1020;
    mem[606] = 'd1020;
    mem[607] = 'd1020;
    mem[608] = 'd1020;
    mem[609] = 'd1020;
    mem[610] = 'd1020;
    mem[611] = 'd1020;
    mem[612] = 'd1020;
    mem[613] = 'd1020;
    mem[614] = 'd1020;
    mem[615] = 'd1020;
    mem[616] = 'd1020;
    mem[617] = 'd1020;
    mem[618] = 'd1020;
    mem[619] = 'd1020;
    mem[620] = 'd1020;
    mem[621] = 'd1020;
    mem[622] = 'd1020;
    mem[623] = 'd1020;
    mem[624] = 'd572;
    mem[625] = 'd804;
    mem[626] = 'd52;
    mem[627] = 'd660;
    mem[628] = 'd52;
    mem[629] = 'd764;
    mem[630] = 'd212;
    mem[631] = 'd868;
    mem[632] = 'd600;
    mem[633] = 'd972;
    mem[634] = 'd840;
    mem[635] = 'd1008;
    mem[636] = 'd852;
    mem[637] = 'd1012;
    mem[638] = 'd864;
    mem[639] = 'd1012;
    mem[640] = 'd880;
    mem[641] = 'd1012;
    mem[642] = 'd888;
    mem[643] = 'd1012;
    mem[644] = 'd892;
    mem[645] = 'd1012;
    mem[646] = 'd892;
    mem[647] = 'd1012;
    mem[648] = 'd888;
    mem[649] = 'd1012;
    mem[650] = 'd876;
    mem[651] = 'd1012;
    mem[652] = 'd864;
    mem[653] = 'd1012;
    mem[654] = 'd848;
    mem[655] = 'd1012;
    mem[656] = 'd836;
    mem[657] = 'd1012;
    mem[658] = 'd648;
    mem[659] = 'd976;
    mem[660] = 'd276;
    mem[661] = 'd880;
    mem[662] = 'd60;
    mem[663] = 'd768;
    mem[664] = 'd84;
    mem[665] = 'd680;
    mem[666] = 'd532;
    mem[667] = 'd792;
    mem[668] = 'd988;
    mem[669] = 'd1004;
    mem[670] = 'd1020;
    mem[671] = 'd1020;
    mem[672] = 'd1020;
    mem[673] = 'd1020;
    mem[674] = 'd1020;
    mem[675] = 'd1020;
    mem[676] = 'd1020;
    mem[677] = 'd1020;
    mem[678] = 'd1020;
    mem[679] = 'd1020;
    mem[680] = 'd1020;
    mem[681] = 'd1020;
    mem[682] = 'd1020;
    mem[683] = 'd1020;
    mem[684] = 'd1020;
    mem[685] = 'd1020;
    mem[686] = 'd1020;
    mem[687] = 'd1020;
    mem[688] = 'd1020;
    mem[689] = 'd1020;
    mem[690] = 'd1020;
    mem[691] = 'd1020;
    mem[692] = 'd1020;
    mem[693] = 'd1020;
    mem[694] = 'd1020;
    mem[695] = 'd1020;
    mem[696] = 'd1020;
    mem[697] = 'd1020;
    mem[698] = 'd1020;
    mem[699] = 'd1020;
    mem[700] = 'd804;
    mem[701] = 'd984;
    mem[702] = 'd660;
    mem[703] = 'd1012;
    mem[704] = 'd764;
    mem[705] = 'd1020;
    mem[706] = 'd868;
    mem[707] = 'd1020;
    mem[708] = 'd972;
    mem[709] = 'd1020;
    mem[710] = 'd1008;
    mem[711] = 'd1020;
    mem[712] = 'd1012;
    mem[713] = 'd1020;
    mem[714] = 'd1012;
    mem[715] = 'd1020;
    mem[716] = 'd1012;
    mem[717] = 'd1020;
    mem[718] = 'd1012;
    mem[719] = 'd1020;
    mem[720] = 'd1012;
    mem[721] = 'd1020;
    mem[722] = 'd1012;
    mem[723] = 'd1020;
    mem[724] = 'd1012;
    mem[725] = 'd1020;
    mem[726] = 'd1012;
    mem[727] = 'd1020;
    mem[728] = 'd1012;
    mem[729] = 'd1020;
    mem[730] = 'd1012;
    mem[731] = 'd1020;
    mem[732] = 'd1012;
    mem[733] = 'd1020;
    mem[734] = 'd976;
    mem[735] = 'd1020;
    mem[736] = 'd880;
    mem[737] = 'd1020;
    mem[738] = 'd768;
    mem[739] = 'd1020;
    mem[740] = 'd680;
    mem[741] = 'd1012;
    mem[742] = 'd792;
    mem[743] = 'd996;
    mem[744] = 'd1004;
    mem[745] = 'd1012;
    mem[746] = 'd1020;
    mem[747] = 'd1020;
    mem[748] = 'd1020;
    mem[749] = 'd1020;
    mem[750] = 'd1020;
    mem[751] = 'd1020;
    mem[752] = 'd1020;
    mem[753] = 'd1020;
    mem[754] = 'd1020;
    mem[755] = 'd1020;
    mem[756] = 'd1020;
    mem[757] = 'd1020;
    mem[758] = 'd1020;
    mem[759] = 'd1020;
    mem[760] = 'd1020;
    mem[761] = 'd1020;
    mem[762] = 'd1020;
    mem[763] = 'd1020;
    mem[764] = 'd1020;
    mem[765] = 'd1020;
    mem[766] = 'd1020;
    mem[767] = 'd1020;
    mem[768] = 'd1020;
    mem[769] = 'd1020;
    mem[770] = 'd1020;
    mem[771] = 'd1020;
    mem[772] = 'd912;
    mem[773] = 'd964;
    mem[774] = 'd296;
    mem[775] = 'd700;
    mem[776] = 'd36;
    mem[777] = 'd696;
    mem[778] = 'd140;
    mem[779] = 'd816;
    mem[780] = 'd520;
    mem[781] = 'd948;
    mem[782] = 'd764;
    mem[783] = 'd1004;
    mem[784] = 'd776;
    mem[785] = 'd1004;
    mem[786] = 'd788;
    mem[787] = 'd1008;
    mem[788] = 'd804;
    mem[789] = 'd1008;
    mem[790] = 'd820;
    mem[791] = 'd1008;
    mem[792] = 'd836;
    mem[793] = 'd1008;
    mem[794] = 'd844;
    mem[795] = 'd1012;
    mem[796] = 'd848;
    mem[797] = 'd1012;
    mem[798] = 'd848;
    mem[799] = 'd1012;
    mem[800] = 'd840;
    mem[801] = 'd1012;
    mem[802] = 'd832;
    mem[803] = 'd1008;
    mem[804] = 'd816;
    mem[805] = 'd1008;
    mem[806] = 'd800;
    mem[807] = 'd1008;
    mem[808] = 'd784;
    mem[809] = 'd1008;
    mem[810] = 'd772;
    mem[811] = 'd1004;
    mem[812] = 'd760;
    mem[813] = 'd1008;
    mem[814] = 'd588;
    mem[815] = 'd964;
    mem[816] = 'd184;
    mem[817] = 'd828;
    mem[818] = 'd36;
    mem[819] = 'd700;
    mem[820] = 'd268;
    mem[821] = 'd688;
    mem[822] = 'd904;
    mem[823] = 'd960;
    mem[824] = 'd1020;
    mem[825] = 'd1020;
    mem[826] = 'd1020;
    mem[827] = 'd1020;
    mem[828] = 'd1020;
    mem[829] = 'd1020;
    mem[830] = 'd1020;
    mem[831] = 'd1020;
    mem[832] = 'd1020;
    mem[833] = 'd1020;
    mem[834] = 'd1020;
    mem[835] = 'd1020;
    mem[836] = 'd1020;
    mem[837] = 'd1020;
    mem[838] = 'd1020;
    mem[839] = 'd1020;
    mem[840] = 'd1020;
    mem[841] = 'd1020;
    mem[842] = 'd1020;
    mem[843] = 'd1020;
    mem[844] = 'd1020;
    mem[845] = 'd1020;
    mem[846] = 'd1020;
    mem[847] = 'd1020;
    mem[848] = 'd964;
    mem[849] = 'd1012;
    mem[850] = 'd700;
    mem[851] = 'd988;
    mem[852] = 'd696;
    mem[853] = 'd1020;
    mem[854] = 'd816;
    mem[855] = 'd1020;
    mem[856] = 'd948;
    mem[857] = 'd1020;
    mem[858] = 'd1004;
    mem[859] = 'd1020;
    mem[860] = 'd1004;
    mem[861] = 'd1020;
    mem[862] = 'd1008;
    mem[863] = 'd1020;
    mem[864] = 'd1008;
    mem[865] = 'd1020;
    mem[866] = 'd1008;
    mem[867] = 'd1020;
    mem[868] = 'd1008;
    mem[869] = 'd1020;
    mem[870] = 'd1012;
    mem[871] = 'd1020;
    mem[872] = 'd1012;
    mem[873] = 'd1020;
    mem[874] = 'd1012;
    mem[875] = 'd1020;
    mem[876] = 'd1012;
    mem[877] = 'd1020;
    mem[878] = 'd1008;
    mem[879] = 'd1020;
    mem[880] = 'd1008;
    mem[881] = 'd1020;
    mem[882] = 'd1008;
    mem[883] = 'd1020;
    mem[884] = 'd1008;
    mem[885] = 'd1020;
    mem[886] = 'd1004;
    mem[887] = 'd1020;
    mem[888] = 'd1008;
    mem[889] = 'd1020;
    mem[890] = 'd964;
    mem[891] = 'd1020;
    mem[892] = 'd828;
    mem[893] = 'd1020;
    mem[894] = 'd700;
    mem[895] = 'd1020;
    mem[896] = 'd688;
    mem[897] = 'd988;
    mem[898] = 'd960;
    mem[899] = 'd1012;
    mem[900] = 'd1020;
    mem[901] = 'd1020;
    mem[902] = 'd1020;
    mem[903] = 'd1020;
    mem[904] = 'd1020;
    mem[905] = 'd1020;
    mem[906] = 'd1020;
    mem[907] = 'd1020;
    mem[908] = 'd1020;
    mem[909] = 'd1020;
    mem[910] = 'd1020;
    mem[911] = 'd1020;
    mem[912] = 'd1020;
    mem[913] = 'd1020;
    mem[914] = 'd1020;
    mem[915] = 'd1020;
    mem[916] = 'd1020;
    mem[917] = 'd1020;
    mem[918] = 'd1020;
    mem[919] = 'd1020;
    mem[920] = 'd1020;
    mem[921] = 'd1020;
    mem[922] = 'd912;
    mem[923] = 'd964;
    mem[924] = 'd188;
    mem[925] = 'd648;
    mem[926] = 'd32;
    mem[927] = 'd708;
    mem[928] = 'd220;
    mem[929] = 'd836;
    mem[930] = 'd632;
    mem[931] = 'd976;
    mem[932] = 'd696;
    mem[933] = 'd1004;
    mem[934] = 'd708;
    mem[935] = 'd1004;
    mem[936] = 'd720;
    mem[937] = 'd1004;
    mem[938] = 'd736;
    mem[939] = 'd1004;
    mem[940] = 'd752;
    mem[941] = 'd1004;
    mem[942] = 'd764;
    mem[943] = 'd1004;
    mem[944] = 'd780;
    mem[945] = 'd1004;
    mem[946] = 'd788;
    mem[947] = 'd1008;
    mem[948] = 'd796;
    mem[949] = 'd1008;
    mem[950] = 'd792;
    mem[951] = 'd1008;
    mem[952] = 'd788;
    mem[953] = 'd1004;
    mem[954] = 'd780;
    mem[955] = 'd1004;
    mem[956] = 'd764;
    mem[957] = 'd1004;
    mem[958] = 'd748;
    mem[959] = 'd1004;
    mem[960] = 'd732;
    mem[961] = 'd1004;
    mem[962] = 'd716;
    mem[963] = 'd1004;
    mem[964] = 'd704;
    mem[965] = 'd1004;
    mem[966] = 'd692;
    mem[967] = 'd1004;
    mem[968] = 'd656;
    mem[969] = 'd980;
    mem[970] = 'd300;
    mem[971] = 'd860;
    mem[972] = 'd32;
    mem[973] = 'd708;
    mem[974] = 'd160;
    mem[975] = 'd644;
    mem[976] = 'd904;
    mem[977] = 'd960;
    mem[978] = 'd1020;
    mem[979] = 'd1020;
    mem[980] = 'd1020;
    mem[981] = 'd1020;
    mem[982] = 'd1020;
    mem[983] = 'd1020;
    mem[984] = 'd1020;
    mem[985] = 'd1020;
    mem[986] = 'd1020;
    mem[987] = 'd1020;
    mem[988] = 'd1020;
    mem[989] = 'd1020;
    mem[990] = 'd1020;
    mem[991] = 'd1020;
    mem[992] = 'd1020;
    mem[993] = 'd1020;
    mem[994] = 'd1020;
    mem[995] = 'd1020;
    mem[996] = 'd1020;
    mem[997] = 'd1020;
    mem[998] = 'd964;
    mem[999] = 'd1008;
    mem[1000] = 'd648;
    mem[1001] = 'd992;
    mem[1002] = 'd708;
    mem[1003] = 'd1020;
    mem[1004] = 'd836;
    mem[1005] = 'd1020;
    mem[1006] = 'd976;
    mem[1007] = 'd1020;
    mem[1008] = 'd1004;
    mem[1009] = 'd1020;
    mem[1010] = 'd1004;
    mem[1011] = 'd1020;
    mem[1012] = 'd1004;
    mem[1013] = 'd1020;
    mem[1014] = 'd1004;
    mem[1015] = 'd1020;
    mem[1016] = 'd1004;
    mem[1017] = 'd1020;
    mem[1018] = 'd1004;
    mem[1019] = 'd1020;
    mem[1020] = 'd1004;
    mem[1021] = 'd1020;
    mem[1022] = 'd1008;
    mem[1023] = 'd1020;
    mem[1024] = 'd1008;
    mem[1025] = 'd1020;
    mem[1026] = 'd1008;
    mem[1027] = 'd1020;
    mem[1028] = 'd1004;
    mem[1029] = 'd1020;
    mem[1030] = 'd1004;
    mem[1031] = 'd1020;
    mem[1032] = 'd1004;
    mem[1033] = 'd1020;
    mem[1034] = 'd1004;
    mem[1035] = 'd1020;
    mem[1036] = 'd1004;
    mem[1037] = 'd1020;
    mem[1038] = 'd1004;
    mem[1039] = 'd1020;
    mem[1040] = 'd1004;
    mem[1041] = 'd1020;
    mem[1042] = 'd1004;
    mem[1043] = 'd1020;
    mem[1044] = 'd980;
    mem[1045] = 'd1020;
    mem[1046] = 'd860;
    mem[1047] = 'd1020;
    mem[1048] = 'd708;
    mem[1049] = 'd1020;
    mem[1050] = 'd644;
    mem[1051] = 'd996;
    mem[1052] = 'd960;
    mem[1053] = 'd1012;
    mem[1054] = 'd1020;
    mem[1055] = 'd1020;
    mem[1056] = 'd1020;
    mem[1057] = 'd1020;
    mem[1058] = 'd1020;
    mem[1059] = 'd1020;
    mem[1060] = 'd1020;
    mem[1061] = 'd1020;
    mem[1062] = 'd1020;
    mem[1063] = 'd1020;
    mem[1064] = 'd1020;
    mem[1065] = 'd1020;
    mem[1066] = 'd1020;
    mem[1067] = 'd1020;
    mem[1068] = 'd1020;
    mem[1069] = 'd1020;
    mem[1070] = 'd1020;
    mem[1071] = 'd1020;
    mem[1072] = 'd964;
    mem[1073] = 'd984;
    mem[1074] = 'd248;
    mem[1075] = 'd660;
    mem[1076] = 'd32;
    mem[1077] = 'd688;
    mem[1078] = 'd232;
    mem[1079] = 'd832;
    mem[1080] = 'd592;
    mem[1081] = 'd960;
    mem[1082] = 'd628;
    mem[1083] = 'd988;
    mem[1084] = 'd640;
    mem[1085] = 'd996;
    mem[1086] = 'd652;
    mem[1087] = 'd1000;
    mem[1088] = 'd664;
    mem[1089] = 'd1000;
    mem[1090] = 'd676;
    mem[1091] = 'd1000;
    mem[1092] = 'd692;
    mem[1093] = 'd1004;
    mem[1094] = 'd708;
    mem[1095] = 'd1004;
    mem[1096] = 'd716;
    mem[1097] = 'd1004;
    mem[1098] = 'd728;
    mem[1099] = 'd1004;
    mem[1100] = 'd732;
    mem[1101] = 'd1004;
    mem[1102] = 'd732;
    mem[1103] = 'd1004;
    mem[1104] = 'd724;
    mem[1105] = 'd1004;
    mem[1106] = 'd716;
    mem[1107] = 'd1004;
    mem[1108] = 'd704;
    mem[1109] = 'd1004;
    mem[1110] = 'd692;
    mem[1111] = 'd1004;
    mem[1112] = 'd676;
    mem[1113] = 'd1000;
    mem[1114] = 'd664;
    mem[1115] = 'd1000;
    mem[1116] = 'd652;
    mem[1117] = 'd1000;
    mem[1118] = 'd640;
    mem[1119] = 'd996;
    mem[1120] = 'd628;
    mem[1121] = 'd988;
    mem[1122] = 'd616;
    mem[1123] = 'd964;
    mem[1124] = 'd300;
    mem[1125] = 'd852;
    mem[1126] = 'd28;
    mem[1127] = 'd692;
    mem[1128] = 'd212;
    mem[1129] = 'd648;
    mem[1130] = 'd948;
    mem[1131] = 'd976;
    mem[1132] = 'd1020;
    mem[1133] = 'd1020;
    mem[1134] = 'd1020;
    mem[1135] = 'd1020;
    mem[1136] = 'd1020;
    mem[1137] = 'd1020;
    mem[1138] = 'd1020;
    mem[1139] = 'd1020;
    mem[1140] = 'd1020;
    mem[1141] = 'd1020;
    mem[1142] = 'd1020;
    mem[1143] = 'd1020;
    mem[1144] = 'd1020;
    mem[1145] = 'd1020;
    mem[1146] = 'd1020;
    mem[1147] = 'd1020;
    mem[1148] = 'd984;
    mem[1149] = 'd1004;
    mem[1150] = 'd660;
    mem[1151] = 'd980;
    mem[1152] = 'd688;
    mem[1153] = 'd1020;
    mem[1154] = 'd832;
    mem[1155] = 'd1020;
    mem[1156] = 'd960;
    mem[1157] = 'd1020;
    mem[1158] = 'd988;
    mem[1159] = 'd1020;
    mem[1160] = 'd996;
    mem[1161] = 'd1020;
    mem[1162] = 'd1000;
    mem[1163] = 'd1020;
    mem[1164] = 'd1000;
    mem[1165] = 'd1020;
    mem[1166] = 'd1000;
    mem[1167] = 'd1020;
    mem[1168] = 'd1004;
    mem[1169] = 'd1020;
    mem[1170] = 'd1004;
    mem[1171] = 'd1020;
    mem[1172] = 'd1004;
    mem[1173] = 'd1020;
    mem[1174] = 'd1004;
    mem[1175] = 'd1020;
    mem[1176] = 'd1004;
    mem[1177] = 'd1020;
    mem[1178] = 'd1004;
    mem[1179] = 'd1020;
    mem[1180] = 'd1004;
    mem[1181] = 'd1020;
    mem[1182] = 'd1004;
    mem[1183] = 'd1020;
    mem[1184] = 'd1004;
    mem[1185] = 'd1020;
    mem[1186] = 'd1004;
    mem[1187] = 'd1020;
    mem[1188] = 'd1000;
    mem[1189] = 'd1020;
    mem[1190] = 'd1000;
    mem[1191] = 'd1020;
    mem[1192] = 'd1000;
    mem[1193] = 'd1020;
    mem[1194] = 'd996;
    mem[1195] = 'd1020;
    mem[1196] = 'd988;
    mem[1197] = 'd1020;
    mem[1198] = 'd964;
    mem[1199] = 'd1020;
    mem[1200] = 'd852;
    mem[1201] = 'd1020;
    mem[1202] = 'd692;
    mem[1203] = 'd1020;
    mem[1204] = 'd648;
    mem[1205] = 'd984;
    mem[1206] = 'd976;
    mem[1207] = 'd1004;
    mem[1208] = 'd1020;
    mem[1209] = 'd1020;
    mem[1210] = 'd1020;
    mem[1211] = 'd1020;
    mem[1212] = 'd1020;
    mem[1213] = 'd1020;
    mem[1214] = 'd1020;
    mem[1215] = 'd1020;
    mem[1216] = 'd1020;
    mem[1217] = 'd1020;
    mem[1218] = 'd1020;
    mem[1219] = 'd1020;
    mem[1220] = 'd1020;
    mem[1221] = 'd1020;
    mem[1222] = 'd1020;
    mem[1223] = 'd1020;
    mem[1224] = 'd452;
    mem[1225] = 'd748;
    mem[1226] = 'd24;
    mem[1227] = 'd656;
    mem[1228] = 'd160;
    mem[1229] = 'd796;
    mem[1230] = 'd524;
    mem[1231] = 'd932;
    mem[1232] = 'd560;
    mem[1233] = 'd964;
    mem[1234] = 'd572;
    mem[1235] = 'd984;
    mem[1236] = 'd584;
    mem[1237] = 'd996;
    mem[1238] = 'd592;
    mem[1239] = 'd996;
    mem[1240] = 'd604;
    mem[1241] = 'd996;
    mem[1242] = 'd616;
    mem[1243] = 'd996;
    mem[1244] = 'd628;
    mem[1245] = 'd996;
    mem[1246] = 'd644;
    mem[1247] = 'd1000;
    mem[1248] = 'd652;
    mem[1249] = 'd1000;
    mem[1250] = 'd660;
    mem[1251] = 'd1000;
    mem[1252] = 'd664;
    mem[1253] = 'd1000;
    mem[1254] = 'd664;
    mem[1255] = 'd1000;
    mem[1256] = 'd660;
    mem[1257] = 'd1000;
    mem[1258] = 'd652;
    mem[1259] = 'd1000;
    mem[1260] = 'd640;
    mem[1261] = 'd1000;
    mem[1262] = 'd628;
    mem[1263] = 'd996;
    mem[1264] = 'd616;
    mem[1265] = 'd996;
    mem[1266] = 'd604;
    mem[1267] = 'd996;
    mem[1268] = 'd592;
    mem[1269] = 'd996;
    mem[1270] = 'd584;
    mem[1271] = 'd996;
    mem[1272] = 'd572;
    mem[1273] = 'd988;
    mem[1274] = 'd560;
    mem[1275] = 'd968;
    mem[1276] = 'd544;
    mem[1277] = 'd936;
    mem[1278] = 'd232;
    mem[1279] = 'd812;
    mem[1280] = 'd24;
    mem[1281] = 'd660;
    mem[1282] = 'd468;
    mem[1283] = 'd752;
    mem[1284] = 'd1020;
    mem[1285] = 'd1020;
    mem[1286] = 'd1020;
    mem[1287] = 'd1020;
    mem[1288] = 'd1020;
    mem[1289] = 'd1020;
    mem[1290] = 'd1020;
    mem[1291] = 'd1020;
    mem[1292] = 'd1020;
    mem[1293] = 'd1020;
    mem[1294] = 'd1020;
    mem[1295] = 'd1020;
    mem[1296] = 'd1020;
    mem[1297] = 'd1020;
    mem[1298] = 'd1020;
    mem[1299] = 'd1020;
    mem[1300] = 'd748;
    mem[1301] = 'd988;
    mem[1302] = 'd656;
    mem[1303] = 'd1020;
    mem[1304] = 'd796;
    mem[1305] = 'd1020;
    mem[1306] = 'd932;
    mem[1307] = 'd1020;
    mem[1308] = 'd964;
    mem[1309] = 'd1020;
    mem[1310] = 'd984;
    mem[1311] = 'd1020;
    mem[1312] = 'd996;
    mem[1313] = 'd1020;
    mem[1314] = 'd996;
    mem[1315] = 'd1020;
    mem[1316] = 'd996;
    mem[1317] = 'd1020;
    mem[1318] = 'd996;
    mem[1319] = 'd1020;
    mem[1320] = 'd996;
    mem[1321] = 'd1020;
    mem[1322] = 'd1000;
    mem[1323] = 'd1020;
    mem[1324] = 'd1000;
    mem[1325] = 'd1020;
    mem[1326] = 'd1000;
    mem[1327] = 'd1020;
    mem[1328] = 'd1000;
    mem[1329] = 'd1020;
    mem[1330] = 'd1000;
    mem[1331] = 'd1020;
    mem[1332] = 'd1000;
    mem[1333] = 'd1020;
    mem[1334] = 'd1000;
    mem[1335] = 'd1020;
    mem[1336] = 'd1000;
    mem[1337] = 'd1020;
    mem[1338] = 'd996;
    mem[1339] = 'd1020;
    mem[1340] = 'd996;
    mem[1341] = 'd1020;
    mem[1342] = 'd996;
    mem[1343] = 'd1020;
    mem[1344] = 'd996;
    mem[1345] = 'd1020;
    mem[1346] = 'd996;
    mem[1347] = 'd1020;
    mem[1348] = 'd988;
    mem[1349] = 'd1020;
    mem[1350] = 'd968;
    mem[1351] = 'd1020;
    mem[1352] = 'd936;
    mem[1353] = 'd1020;
    mem[1354] = 'd812;
    mem[1355] = 'd1020;
    mem[1356] = 'd660;
    mem[1357] = 'd1020;
    mem[1358] = 'd752;
    mem[1359] = 'd984;
    mem[1360] = 'd1020;
    mem[1361] = 'd1020;
    mem[1362] = 'd1020;
    mem[1363] = 'd1020;
    mem[1364] = 'd1020;
    mem[1365] = 'd1020;
    mem[1366] = 'd1020;
    mem[1367] = 'd1020;
    mem[1368] = 'd1020;
    mem[1369] = 'd1020;
    mem[1370] = 'd1020;
    mem[1371] = 'd1020;
    mem[1372] = 'd1020;
    mem[1373] = 'd1020;
    mem[1374] = 'd840;
    mem[1375] = 'd924;
    mem[1376] = 'd32;
    mem[1377] = 'd608;
    mem[1378] = 'd76;
    mem[1379] = 'd736;
    mem[1380] = 'd436;
    mem[1381] = 'd896;
    mem[1382] = 'd496;
    mem[1383] = 'd936;
    mem[1384] = 'd508;
    mem[1385] = 'd956;
    mem[1386] = 'd516;
    mem[1387] = 'd976;
    mem[1388] = 'd528;
    mem[1389] = 'd992;
    mem[1390] = 'd536;
    mem[1391] = 'd992;
    mem[1392] = 'd544;
    mem[1393] = 'd996;
    mem[1394] = 'd556;
    mem[1395] = 'd996;
    mem[1396] = 'd568;
    mem[1397] = 'd996;
    mem[1398] = 'd576;
    mem[1399] = 'd996;
    mem[1400] = 'd584;
    mem[1401] = 'd996;
    mem[1402] = 'd592;
    mem[1403] = 'd996;
    mem[1404] = 'd596;
    mem[1405] = 'd996;
    mem[1406] = 'd596;
    mem[1407] = 'd996;
    mem[1408] = 'd592;
    mem[1409] = 'd996;
    mem[1410] = 'd584;
    mem[1411] = 'd996;
    mem[1412] = 'd576;
    mem[1413] = 'd996;
    mem[1414] = 'd564;
    mem[1415] = 'd996;
    mem[1416] = 'd556;
    mem[1417] = 'd996;
    mem[1418] = 'd544;
    mem[1419] = 'd996;
    mem[1420] = 'd532;
    mem[1421] = 'd992;
    mem[1422] = 'd524;
    mem[1423] = 'd992;
    mem[1424] = 'd516;
    mem[1425] = 'd976;
    mem[1426] = 'd508;
    mem[1427] = 'd956;
    mem[1428] = 'd496;
    mem[1429] = 'd936;
    mem[1430] = 'd460;
    mem[1431] = 'd900;
    mem[1432] = 'd116;
    mem[1433] = 'd748;
    mem[1434] = 'd28;
    mem[1435] = 'd604;
    mem[1436] = 'd828;
    mem[1437] = 'd912;
    mem[1438] = 'd1020;
    mem[1439] = 'd1020;
    mem[1440] = 'd1020;
    mem[1441] = 'd1020;
    mem[1442] = 'd1020;
    mem[1443] = 'd1020;
    mem[1444] = 'd1020;
    mem[1445] = 'd1020;
    mem[1446] = 'd1020;
    mem[1447] = 'd1020;
    mem[1448] = 'd1020;
    mem[1449] = 'd1020;
    mem[1450] = 'd924;
    mem[1451] = 'd996;
    mem[1452] = 'd608;
    mem[1453] = 'd1008;
    mem[1454] = 'd736;
    mem[1455] = 'd1020;
    mem[1456] = 'd896;
    mem[1457] = 'd1020;
    mem[1458] = 'd936;
    mem[1459] = 'd1020;
    mem[1460] = 'd956;
    mem[1461] = 'd1020;
    mem[1462] = 'd976;
    mem[1463] = 'd1020;
    mem[1464] = 'd992;
    mem[1465] = 'd1020;
    mem[1466] = 'd992;
    mem[1467] = 'd1020;
    mem[1468] = 'd996;
    mem[1469] = 'd1020;
    mem[1470] = 'd996;
    mem[1471] = 'd1020;
    mem[1472] = 'd996;
    mem[1473] = 'd1020;
    mem[1474] = 'd996;
    mem[1475] = 'd1020;
    mem[1476] = 'd996;
    mem[1477] = 'd1020;
    mem[1478] = 'd996;
    mem[1479] = 'd1020;
    mem[1480] = 'd996;
    mem[1481] = 'd1020;
    mem[1482] = 'd996;
    mem[1483] = 'd1020;
    mem[1484] = 'd996;
    mem[1485] = 'd1020;
    mem[1486] = 'd996;
    mem[1487] = 'd1020;
    mem[1488] = 'd996;
    mem[1489] = 'd1020;
    mem[1490] = 'd996;
    mem[1491] = 'd1020;
    mem[1492] = 'd996;
    mem[1493] = 'd1020;
    mem[1494] = 'd996;
    mem[1495] = 'd1020;
    mem[1496] = 'd992;
    mem[1497] = 'd1020;
    mem[1498] = 'd992;
    mem[1499] = 'd1020;
    mem[1500] = 'd976;
    mem[1501] = 'd1020;
    mem[1502] = 'd956;
    mem[1503] = 'd1020;
    mem[1504] = 'd936;
    mem[1505] = 'd1020;
    mem[1506] = 'd900;
    mem[1507] = 'd1020;
    mem[1508] = 'd748;
    mem[1509] = 'd1020;
    mem[1510] = 'd604;
    mem[1511] = 'd1012;
    mem[1512] = 'd912;
    mem[1513] = 'd988;
    mem[1514] = 'd1020;
    mem[1515] = 'd1020;
    mem[1516] = 'd1020;
    mem[1517] = 'd1020;
    mem[1518] = 'd1020;
    mem[1519] = 'd1020;
    mem[1520] = 'd1020;
    mem[1521] = 'd1020;
    mem[1522] = 'd1020;
    mem[1523] = 'd1020;
    mem[1524] = 'd1012;
    mem[1525] = 'd1016;
    mem[1526] = 'd304;
    mem[1527] = 'd668;
    mem[1528] = 'd32;
    mem[1529] = 'd668;
    mem[1530] = 'd284;
    mem[1531] = 'd824;
    mem[1532] = 'd428;
    mem[1533] = 'd900;
    mem[1534] = 'd440;
    mem[1535] = 'd924;
    mem[1536] = 'd452;
    mem[1537] = 'd948;
    mem[1538] = 'd456;
    mem[1539] = 'd964;
    mem[1540] = 'd464;
    mem[1541] = 'd976;
    mem[1542] = 'd476;
    mem[1543] = 'd988;
    mem[1544] = 'd484;
    mem[1545] = 'd988;
    mem[1546] = 'd492;
    mem[1547] = 'd988;
    mem[1548] = 'd504;
    mem[1549] = 'd992;
    mem[1550] = 'd512;
    mem[1551] = 'd992;
    mem[1552] = 'd520;
    mem[1553] = 'd992;
    mem[1554] = 'd524;
    mem[1555] = 'd992;
    mem[1556] = 'd528;
    mem[1557] = 'd992;
    mem[1558] = 'd528;
    mem[1559] = 'd992;
    mem[1560] = 'd524;
    mem[1561] = 'd992;
    mem[1562] = 'd520;
    mem[1563] = 'd992;
    mem[1564] = 'd508;
    mem[1565] = 'd992;
    mem[1566] = 'd504;
    mem[1567] = 'd992;
    mem[1568] = 'd492;
    mem[1569] = 'd988;
    mem[1570] = 'd484;
    mem[1571] = 'd988;
    mem[1572] = 'd476;
    mem[1573] = 'd988;
    mem[1574] = 'd464;
    mem[1575] = 'd976;
    mem[1576] = 'd460;
    mem[1577] = 'd964;
    mem[1578] = 'd448;
    mem[1579] = 'd948;
    mem[1580] = 'd440;
    mem[1581] = 'd928;
    mem[1582] = 'd428;
    mem[1583] = 'd900;
    mem[1584] = 'd336;
    mem[1585] = 'd844;
    mem[1586] = 'd40;
    mem[1587] = 'd672;
    mem[1588] = 'd256;
    mem[1589] = 'd644;
    mem[1590] = 'd1020;
    mem[1591] = 'd1020;
    mem[1592] = 'd1020;
    mem[1593] = 'd1020;
    mem[1594] = 'd1020;
    mem[1595] = 'd1020;
    mem[1596] = 'd1020;
    mem[1597] = 'd1020;
    mem[1598] = 'd1020;
    mem[1599] = 'd1020;
    mem[1600] = 'd1016;
    mem[1601] = 'd1016;
    mem[1602] = 'd668;
    mem[1603] = 'd972;
    mem[1604] = 'd668;
    mem[1605] = 'd1020;
    mem[1606] = 'd824;
    mem[1607] = 'd1020;
    mem[1608] = 'd900;
    mem[1609] = 'd1020;
    mem[1610] = 'd924;
    mem[1611] = 'd1020;
    mem[1612] = 'd948;
    mem[1613] = 'd1020;
    mem[1614] = 'd964;
    mem[1615] = 'd1020;
    mem[1616] = 'd976;
    mem[1617] = 'd1020;
    mem[1618] = 'd988;
    mem[1619] = 'd1020;
    mem[1620] = 'd988;
    mem[1621] = 'd1020;
    mem[1622] = 'd988;
    mem[1623] = 'd1020;
    mem[1624] = 'd992;
    mem[1625] = 'd1020;
    mem[1626] = 'd992;
    mem[1627] = 'd1020;
    mem[1628] = 'd992;
    mem[1629] = 'd1020;
    mem[1630] = 'd992;
    mem[1631] = 'd1020;
    mem[1632] = 'd992;
    mem[1633] = 'd1020;
    mem[1634] = 'd992;
    mem[1635] = 'd1020;
    mem[1636] = 'd992;
    mem[1637] = 'd1020;
    mem[1638] = 'd992;
    mem[1639] = 'd1020;
    mem[1640] = 'd992;
    mem[1641] = 'd1020;
    mem[1642] = 'd992;
    mem[1643] = 'd1020;
    mem[1644] = 'd988;
    mem[1645] = 'd1020;
    mem[1646] = 'd988;
    mem[1647] = 'd1020;
    mem[1648] = 'd988;
    mem[1649] = 'd1020;
    mem[1650] = 'd976;
    mem[1651] = 'd1020;
    mem[1652] = 'd964;
    mem[1653] = 'd1020;
    mem[1654] = 'd948;
    mem[1655] = 'd1020;
    mem[1656] = 'd928;
    mem[1657] = 'd1020;
    mem[1658] = 'd900;
    mem[1659] = 'd1020;
    mem[1660] = 'd844;
    mem[1661] = 'd1020;
    mem[1662] = 'd672;
    mem[1663] = 'd1020;
    mem[1664] = 'd644;
    mem[1665] = 'd972;
    mem[1666] = 'd1020;
    mem[1667] = 'd1020;
    mem[1668] = 'd1020;
    mem[1669] = 'd1020;
    mem[1670] = 'd1020;
    mem[1671] = 'd1020;
    mem[1672] = 'd1020;
    mem[1673] = 'd1020;
    mem[1674] = 'd1020;
    mem[1675] = 'd1020;
    mem[1676] = 'd788;
    mem[1677] = 'd892;
    mem[1678] = 'd24;
    mem[1679] = 'd584;
    mem[1680] = 'd108;
    mem[1681] = 'd700;
    mem[1682] = 'd344;
    mem[1683] = 'd804;
    mem[1684] = 'd356;
    mem[1685] = 'd824;
    mem[1686] = 'd364;
    mem[1687] = 'd840;
    mem[1688] = 'd372;
    mem[1689] = 'd860;
    mem[1690] = 'd388;
    mem[1691] = 'd888;
    mem[1692] = 'd396;
    mem[1693] = 'd912;
    mem[1694] = 'd408;
    mem[1695] = 'd952;
    mem[1696] = 'd424;
    mem[1697] = 'd988;
    mem[1698] = 'd436;
    mem[1699] = 'd992;
    mem[1700] = 'd436;
    mem[1701] = 'd988;
    mem[1702] = 'd448;
    mem[1703] = 'd988;
    mem[1704] = 'd456;
    mem[1705] = 'd988;
    mem[1706] = 'd456;
    mem[1707] = 'd988;
    mem[1708] = 'd460;
    mem[1709] = 'd988;
    mem[1710] = 'd460;
    mem[1711] = 'd988;
    mem[1712] = 'd460;
    mem[1713] = 'd988;
    mem[1714] = 'd456;
    mem[1715] = 'd988;
    mem[1716] = 'd444;
    mem[1717] = 'd988;
    mem[1718] = 'd436;
    mem[1719] = 'd992;
    mem[1720] = 'd432;
    mem[1721] = 'd992;
    mem[1722] = 'd424;
    mem[1723] = 'd980;
    mem[1724] = 'd404;
    mem[1725] = 'd944;
    mem[1726] = 'd392;
    mem[1727] = 'd908;
    mem[1728] = 'd380;
    mem[1729] = 'd884;
    mem[1730] = 'd376;
    mem[1731] = 'd860;
    mem[1732] = 'd368;
    mem[1733] = 'd844;
    mem[1734] = 'd356;
    mem[1735] = 'd828;
    mem[1736] = 'd348;
    mem[1737] = 'd812;
    mem[1738] = 'd148;
    mem[1739] = 'd728;
    mem[1740] = 'd16;
    mem[1741] = 'd584;
    mem[1742] = 'd760;
    mem[1743] = 'd872;
    mem[1744] = 'd1020;
    mem[1745] = 'd1020;
    mem[1746] = 'd1020;
    mem[1747] = 'd1020;
    mem[1748] = 'd1020;
    mem[1749] = 'd1020;
    mem[1750] = 'd1020;
    mem[1751] = 'd1020;
    mem[1752] = 'd892;
    mem[1753] = 'd984;
    mem[1754] = 'd584;
    mem[1755] = 'd1000;
    mem[1756] = 'd700;
    mem[1757] = 'd968;
    mem[1758] = 'd804;
    mem[1759] = 'd948;
    mem[1760] = 'd824;
    mem[1761] = 'd940;
    mem[1762] = 'd840;
    mem[1763] = 'd932;
    mem[1764] = 'd860;
    mem[1765] = 'd936;
    mem[1766] = 'd888;
    mem[1767] = 'd944;
    mem[1768] = 'd912;
    mem[1769] = 'd956;
    mem[1770] = 'd952;
    mem[1771] = 'd980;
    mem[1772] = 'd988;
    mem[1773] = 'd1012;
    mem[1774] = 'd992;
    mem[1775] = 'd1020;
    mem[1776] = 'd988;
    mem[1777] = 'd1020;
    mem[1778] = 'd988;
    mem[1779] = 'd1020;
    mem[1780] = 'd988;
    mem[1781] = 'd1020;
    mem[1782] = 'd988;
    mem[1783] = 'd1020;
    mem[1784] = 'd988;
    mem[1785] = 'd1020;
    mem[1786] = 'd988;
    mem[1787] = 'd1020;
    mem[1788] = 'd988;
    mem[1789] = 'd1020;
    mem[1790] = 'd988;
    mem[1791] = 'd1020;
    mem[1792] = 'd988;
    mem[1793] = 'd1020;
    mem[1794] = 'd992;
    mem[1795] = 'd1020;
    mem[1796] = 'd992;
    mem[1797] = 'd1020;
    mem[1798] = 'd980;
    mem[1799] = 'd1008;
    mem[1800] = 'd944;
    mem[1801] = 'd976;
    mem[1802] = 'd908;
    mem[1803] = 'd956;
    mem[1804] = 'd884;
    mem[1805] = 'd940;
    mem[1806] = 'd860;
    mem[1807] = 'd932;
    mem[1808] = 'd844;
    mem[1809] = 'd936;
    mem[1810] = 'd828;
    mem[1811] = 'd940;
    mem[1812] = 'd812;
    mem[1813] = 'd952;
    mem[1814] = 'd728;
    mem[1815] = 'd988;
    mem[1816] = 'd584;
    mem[1817] = 'd1004;
    mem[1818] = 'd872;
    mem[1819] = 'd976;
    mem[1820] = 'd1020;
    mem[1821] = 'd1020;
    mem[1822] = 'd1020;
    mem[1823] = 'd1020;
    mem[1824] = 'd1020;
    mem[1825] = 'd1020;
    mem[1826] = 'd1020;
    mem[1827] = 'd1020;
    mem[1828] = 'd352;
    mem[1829] = 'd676;
    mem[1830] = 'd52;
    mem[1831] = 'd460;
    mem[1832] = 'd132;
    mem[1833] = 'd168;
    mem[1834] = 'd152;
    mem[1835] = 'd168;
    mem[1836] = 'd152;
    mem[1837] = 'd168;
    mem[1838] = 'd148;
    mem[1839] = 'd160;
    mem[1840] = 'd140;
    mem[1841] = 'd152;
    mem[1842] = 'd144;
    mem[1843] = 'd160;
    mem[1844] = 'd152;
    mem[1845] = 'd176;
    mem[1846] = 'd172;
    mem[1847] = 'd220;
    mem[1848] = 'd204;
    mem[1849] = 'd304;
    mem[1850] = 'd248;
    mem[1851] = 'd428;
    mem[1852] = 'd308;
    mem[1853] = 'd628;
    mem[1854] = 'd340;
    mem[1855] = 'd820;
    mem[1856] = 'd392;
    mem[1857] = 'd980;
    mem[1858] = 'd396;
    mem[1859] = 'd988;
    mem[1860] = 'd396;
    mem[1861] = 'd984;
    mem[1862] = 'd396;
    mem[1863] = 'd988;
    mem[1864] = 'd396;
    mem[1865] = 'd988;
    mem[1866] = 'd380;
    mem[1867] = 'd944;
    mem[1868] = 'd336;
    mem[1869] = 'd788;
    mem[1870] = 'd296;
    mem[1871] = 'd596;
    mem[1872] = 'd244;
    mem[1873] = 'd408;
    mem[1874] = 'd200;
    mem[1875] = 'd288;
    mem[1876] = 'd172;
    mem[1877] = 'd212;
    mem[1878] = 'd152;
    mem[1879] = 'd172;
    mem[1880] = 'd144;
    mem[1881] = 'd164;
    mem[1882] = 'd144;
    mem[1883] = 'd156;
    mem[1884] = 'd156;
    mem[1885] = 'd168;
    mem[1886] = 'd156;
    mem[1887] = 'd172;
    mem[1888] = 'd152;
    mem[1889] = 'd172;
    mem[1890] = 'd132;
    mem[1891] = 'd168;
    mem[1892] = 'd44;
    mem[1893] = 'd540;
    mem[1894] = 'd332;
    mem[1895] = 'd668;
    mem[1896] = 'd1020;
    mem[1897] = 'd1020;
    mem[1898] = 'd1020;
    mem[1899] = 'd1020;
    mem[1900] = 'd1020;
    mem[1901] = 'd1020;
    mem[1902] = 'd1020;
    mem[1903] = 'd1020;
    mem[1904] = 'd676;
    mem[1905] = 'd952;
    mem[1906] = 'd460;
    mem[1907] = 'd732;
    mem[1908] = 'd168;
    mem[1909] = 'd184;
    mem[1910] = 'd168;
    mem[1911] = 'd172;
    mem[1912] = 'd168;
    mem[1913] = 'd168;
    mem[1914] = 'd160;
    mem[1915] = 'd160;
    mem[1916] = 'd152;
    mem[1917] = 'd156;
    mem[1918] = 'd160;
    mem[1919] = 'd160;
    mem[1920] = 'd176;
    mem[1921] = 'd176;
    mem[1922] = 'd220;
    mem[1923] = 'd220;
    mem[1924] = 'd304;
    mem[1925] = 'd308;
    mem[1926] = 'd428;
    mem[1927] = 'd436;
    mem[1928] = 'd628;
    mem[1929] = 'd636;
    mem[1930] = 'd820;
    mem[1931] = 'd840;
    mem[1932] = 'd980;
    mem[1933] = 'd1004;
    mem[1934] = 'd988;
    mem[1935] = 'd1020;
    mem[1936] = 'd984;
    mem[1937] = 'd1020;
    mem[1938] = 'd988;
    mem[1939] = 'd1020;
    mem[1940] = 'd988;
    mem[1941] = 'd1020;
    mem[1942] = 'd944;
    mem[1943] = 'd972;
    mem[1944] = 'd788;
    mem[1945] = 'd804;
    mem[1946] = 'd596;
    mem[1947] = 'd608;
    mem[1948] = 'd408;
    mem[1949] = 'd412;
    mem[1950] = 'd288;
    mem[1951] = 'd296;
    mem[1952] = 'd212;
    mem[1953] = 'd216;
    mem[1954] = 'd172;
    mem[1955] = 'd176;
    mem[1956] = 'd164;
    mem[1957] = 'd160;
    mem[1958] = 'd156;
    mem[1959] = 'd160;
    mem[1960] = 'd168;
    mem[1961] = 'd172;
    mem[1962] = 'd172;
    mem[1963] = 'd176;
    mem[1964] = 'd172;
    mem[1965] = 'd180;
    mem[1966] = 'd168;
    mem[1967] = 'd184;
    mem[1968] = 'd540;
    mem[1969] = 'd860;
    mem[1970] = 'd668;
    mem[1971] = 'd956;
    mem[1972] = 'd1020;
    mem[1973] = 'd1020;
    mem[1974] = 'd1020;
    mem[1975] = 'd1020;
    mem[1976] = 'd1020;
    mem[1977] = 'd1020;
    mem[1978] = 'd936;
    mem[1979] = 'd976;
    mem[1980] = 'd76;
    mem[1981] = 'd564;
    mem[1982] = 'd56;
    mem[1983] = 'd488;
    mem[1984] = 'd88;
    mem[1985] = 'd84;
    mem[1986] = 'd88;
    mem[1987] = 'd88;
    mem[1988] = 'd160;
    mem[1989] = 'd164;
    mem[1990] = 'd432;
    mem[1991] = 'd440;
    mem[1992] = 'd532;
    mem[1993] = 'd544;
    mem[1994] = 'd580;
    mem[1995] = 'd596;
    mem[1996] = 'd596;
    mem[1997] = 'd608;
    mem[1998] = 'd576;
    mem[1999] = 'd588;
    mem[2000] = 'd512;
    mem[2001] = 'd524;
    mem[2002] = 'd412;
    mem[2003] = 'd424;
    mem[2004] = 'd264;
    mem[2005] = 'd268;
    mem[2006] = 'd152;
    mem[2007] = 'd152;
    mem[2008] = 'd192;
    mem[2009] = 'd268;
    mem[2010] = 'd268;
    mem[2011] = 'd508;
    mem[2012] = 'd296;
    mem[2013] = 'd612;
    mem[2014] = 'd284;
    mem[2015] = 'd596;
    mem[2016] = 'd248;
    mem[2017] = 'd472;
    mem[2018] = 'd176;
    mem[2019] = 'd248;
    mem[2020] = 'd180;
    mem[2021] = 'd184;
    mem[2022] = 'd288;
    mem[2023] = 'd292;
    mem[2024] = 'd412;
    mem[2025] = 'd420;
    mem[2026] = 'd488;
    mem[2027] = 'd500;
    mem[2028] = 'd540;
    mem[2029] = 'd548;
    mem[2030] = 'd548;
    mem[2031] = 'd560;
    mem[2032] = 'd528;
    mem[2033] = 'd536;
    mem[2034] = 'd468;
    mem[2035] = 'd480;
    mem[2036] = 'd340;
    mem[2037] = 'd348;
    mem[2038] = 'd116;
    mem[2039] = 'd116;
    mem[2040] = 'd88;
    mem[2041] = 'd88;
    mem[2042] = 'd92;
    mem[2043] = 'd100;
    mem[2044] = 'd44;
    mem[2045] = 'd524;
    mem[2046] = 'd28;
    mem[2047] = 'd536;
    mem[2048] = 'd952;
    mem[2049] = 'd984;
    mem[2050] = 'd1020;
    mem[2051] = 'd1020;
    mem[2052] = 'd1020;
    mem[2053] = 'd1020;
    mem[2054] = 'd976;
    mem[2055] = 'd1000;
    mem[2056] = 'd564;
    mem[2057] = 'd940;
    mem[2058] = 'd488;
    mem[2059] = 'd744;
    mem[2060] = 'd84;
    mem[2061] = 'd84;
    mem[2062] = 'd88;
    mem[2063] = 'd88;
    mem[2064] = 'd164;
    mem[2065] = 'd164;
    mem[2066] = 'd440;
    mem[2067] = 'd432;
    mem[2068] = 'd544;
    mem[2069] = 'd536;
    mem[2070] = 'd596;
    mem[2071] = 'd584;
    mem[2072] = 'd608;
    mem[2073] = 'd600;
    mem[2074] = 'd588;
    mem[2075] = 'd576;
    mem[2076] = 'd524;
    mem[2077] = 'd516;
    mem[2078] = 'd424;
    mem[2079] = 'd416;
    mem[2080] = 'd268;
    mem[2081] = 'd264;
    mem[2082] = 'd152;
    mem[2083] = 'd152;
    mem[2084] = 'd268;
    mem[2085] = 'd272;
    mem[2086] = 'd508;
    mem[2087] = 'd516;
    mem[2088] = 'd612;
    mem[2089] = 'd620;
    mem[2090] = 'd596;
    mem[2091] = 'd604;
    mem[2092] = 'd472;
    mem[2093] = 'd480;
    mem[2094] = 'd248;
    mem[2095] = 'd252;
    mem[2096] = 'd184;
    mem[2097] = 'd184;
    mem[2098] = 'd292;
    mem[2099] = 'd288;
    mem[2100] = 'd420;
    mem[2101] = 'd416;
    mem[2102] = 'd500;
    mem[2103] = 'd492;
    mem[2104] = 'd548;
    mem[2105] = 'd540;
    mem[2106] = 'd560;
    mem[2107] = 'd548;
    mem[2108] = 'd536;
    mem[2109] = 'd528;
    mem[2110] = 'd480;
    mem[2111] = 'd468;
    mem[2112] = 'd348;
    mem[2113] = 'd340;
    mem[2114] = 'd116;
    mem[2115] = 'd116;
    mem[2116] = 'd88;
    mem[2117] = 'd88;
    mem[2118] = 'd100;
    mem[2119] = 'd100;
    mem[2120] = 'd524;
    mem[2121] = 'd796;
    mem[2122] = 'd536;
    mem[2123] = 'd932;
    mem[2124] = 'd984;
    mem[2125] = 'd1004;
    mem[2126] = 'd1020;
    mem[2127] = 'd1020;
    mem[2128] = 'd1020;
    mem[2129] = 'd1020;
    mem[2130] = 'd720;
    mem[2131] = 'd852;
    mem[2132] = 'd16;
    mem[2133] = 'd552;
    mem[2134] = 'd52;
    mem[2135] = 'd632;
    mem[2136] = 'd92;
    mem[2137] = 'd152;
    mem[2138] = 'd84;
    mem[2139] = 'd84;
    mem[2140] = 'd328;
    mem[2141] = 'd332;
    mem[2142] = 'd452;
    mem[2143] = 'd464;
    mem[2144] = 'd508;
    mem[2145] = 'd520;
    mem[2146] = 'd532;
    mem[2147] = 'd544;
    mem[2148] = 'd536;
    mem[2149] = 'd552;
    mem[2150] = 'd540;
    mem[2151] = 'd552;
    mem[2152] = 'd536;
    mem[2153] = 'd548;
    mem[2154] = 'd540;
    mem[2155] = 'd556;
    mem[2156] = 'd564;
    mem[2157] = 'd576;
    mem[2158] = 'd520;
    mem[2159] = 'd532;
    mem[2160] = 'd196;
    mem[2161] = 'd200;
    mem[2162] = 'd100;
    mem[2163] = 'd104;
    mem[2164] = 'd144;
    mem[2165] = 'd144;
    mem[2166] = 'd128;
    mem[2167] = 'd128;
    mem[2168] = 'd100;
    mem[2169] = 'd100;
    mem[2170] = 'd248;
    mem[2171] = 'd252;
    mem[2172] = 'd464;
    mem[2173] = 'd476;
    mem[2174] = 'd480;
    mem[2175] = 'd492;
    mem[2176] = 'd460;
    mem[2177] = 'd472;
    mem[2178] = 'd456;
    mem[2179] = 'd464;
    mem[2180] = 'd452;
    mem[2181] = 'd460;
    mem[2182] = 'd440;
    mem[2183] = 'd452;
    mem[2184] = 'd420;
    mem[2185] = 'd432;
    mem[2186] = 'd388;
    mem[2187] = 'd396;
    mem[2188] = 'd328;
    mem[2189] = 'd336;
    mem[2190] = 'd208;
    mem[2191] = 'd212;
    mem[2192] = 'd84;
    mem[2193] = 'd84;
    mem[2194] = 'd84;
    mem[2195] = 'd212;
    mem[2196] = 'd40;
    mem[2197] = 'd596;
    mem[2198] = 'd12;
    mem[2199] = 'd556;
    mem[2200] = 'd652;
    mem[2201] = 'd816;
    mem[2202] = 'd1020;
    mem[2203] = 'd1020;
    mem[2204] = 'd1020;
    mem[2205] = 'd1020;
    mem[2206] = 'd852;
    mem[2207] = 'd972;
    mem[2208] = 'd552;
    mem[2209] = 'd948;
    mem[2210] = 'd632;
    mem[2211] = 'd952;
    mem[2212] = 'd152;
    mem[2213] = 'd184;
    mem[2214] = 'd84;
    mem[2215] = 'd84;
    mem[2216] = 'd332;
    mem[2217] = 'd328;
    mem[2218] = 'd464;
    mem[2219] = 'd452;
    mem[2220] = 'd520;
    mem[2221] = 'd512;
    mem[2222] = 'd544;
    mem[2223] = 'd536;
    mem[2224] = 'd552;
    mem[2225] = 'd540;
    mem[2226] = 'd552;
    mem[2227] = 'd540;
    mem[2228] = 'd548;
    mem[2229] = 'd540;
    mem[2230] = 'd556;
    mem[2231] = 'd544;
    mem[2232] = 'd576;
    mem[2233] = 'd564;
    mem[2234] = 'd532;
    mem[2235] = 'd520;
    mem[2236] = 'd200;
    mem[2237] = 'd196;
    mem[2238] = 'd104;
    mem[2239] = 'd100;
    mem[2240] = 'd144;
    mem[2241] = 'd144;
    mem[2242] = 'd128;
    mem[2243] = 'd128;
    mem[2244] = 'd100;
    mem[2245] = 'd100;
    mem[2246] = 'd252;
    mem[2247] = 'd248;
    mem[2248] = 'd476;
    mem[2249] = 'd464;
    mem[2250] = 'd492;
    mem[2251] = 'd484;
    mem[2252] = 'd472;
    mem[2253] = 'd460;
    mem[2254] = 'd464;
    mem[2255] = 'd456;
    mem[2256] = 'd460;
    mem[2257] = 'd452;
    mem[2258] = 'd452;
    mem[2259] = 'd444;
    mem[2260] = 'd432;
    mem[2261] = 'd424;
    mem[2262] = 'd396;
    mem[2263] = 'd388;
    mem[2264] = 'd336;
    mem[2265] = 'd332;
    mem[2266] = 'd212;
    mem[2267] = 'd208;
    mem[2268] = 'd84;
    mem[2269] = 'd84;
    mem[2270] = 'd212;
    mem[2271] = 'd280;
    mem[2272] = 'd596;
    mem[2273] = 'd896;
    mem[2274] = 'd556;
    mem[2275] = 'd932;
    mem[2276] = 'd816;
    mem[2277] = 'd960;
    mem[2278] = 'd1020;
    mem[2279] = 'd1020;
    mem[2280] = 'd1020;
    mem[2281] = 'd1020;
    mem[2282] = 'd464;
    mem[2283] = 'd716;
    mem[2284] = 'd20;
    mem[2285] = 'd572;
    mem[2286] = 'd72;
    mem[2287] = 'd640;
    mem[2288] = 'd96;
    mem[2289] = 'd384;
    mem[2290] = 'd92;
    mem[2291] = 'd88;
    mem[2292] = 'd212;
    mem[2293] = 'd216;
    mem[2294] = 'd252;
    mem[2295] = 'd256;
    mem[2296] = 'd260;
    mem[2297] = 'd268;
    mem[2298] = 'd272;
    mem[2299] = 'd280;
    mem[2300] = 'd280;
    mem[2301] = 'd292;
    mem[2302] = 'd280;
    mem[2303] = 'd288;
    mem[2304] = 'd264;
    mem[2305] = 'd268;
    mem[2306] = 'd244;
    mem[2307] = 'd252;
    mem[2308] = 'd232;
    mem[2309] = 'd236;
    mem[2310] = 'd216;
    mem[2311] = 'd224;
    mem[2312] = 'd144;
    mem[2313] = 'd148;
    mem[2314] = 'd84;
    mem[2315] = 'd84;
    mem[2316] = 'd76;
    mem[2317] = 'd264;
    mem[2318] = 'd76;
    mem[2319] = 'd188;
    mem[2320] = 'd84;
    mem[2321] = 'd84;
    mem[2322] = 'd148;
    mem[2323] = 'd152;
    mem[2324] = 'd180;
    mem[2325] = 'd184;
    mem[2326] = 'd180;
    mem[2327] = 'd188;
    mem[2328] = 'd184;
    mem[2329] = 'd188;
    mem[2330] = 'd192;
    mem[2331] = 'd196;
    mem[2332] = 'd196;
    mem[2333] = 'd200;
    mem[2334] = 'd184;
    mem[2335] = 'd188;
    mem[2336] = 'd168;
    mem[2337] = 'd172;
    mem[2338] = 'd148;
    mem[2339] = 'd156;
    mem[2340] = 'd136;
    mem[2341] = 'd140;
    mem[2342] = 'd104;
    mem[2343] = 'd104;
    mem[2344] = 'd92;
    mem[2345] = 'd88;
    mem[2346] = 'd68;
    mem[2347] = 'd420;
    mem[2348] = 'd56;
    mem[2349] = 'd612;
    mem[2350] = 'd20;
    mem[2351] = 'd572;
    mem[2352] = 'd420;
    mem[2353] = 'd692;
    mem[2354] = 'd1020;
    mem[2355] = 'd1020;
    mem[2356] = 'd1020;
    mem[2357] = 'd1020;
    mem[2358] = 'd716;
    mem[2359] = 'd940;
    mem[2360] = 'd572;
    mem[2361] = 'd956;
    mem[2362] = 'd640;
    mem[2363] = 'd948;
    mem[2364] = 'd384;
    mem[2365] = 'd524;
    mem[2366] = 'd88;
    mem[2367] = 'd88;
    mem[2368] = 'd216;
    mem[2369] = 'd212;
    mem[2370] = 'd256;
    mem[2371] = 'd252;
    mem[2372] = 'd268;
    mem[2373] = 'd264;
    mem[2374] = 'd280;
    mem[2375] = 'd276;
    mem[2376] = 'd292;
    mem[2377] = 'd284;
    mem[2378] = 'd288;
    mem[2379] = 'd280;
    mem[2380] = 'd268;
    mem[2381] = 'd264;
    mem[2382] = 'd252;
    mem[2383] = 'd244;
    mem[2384] = 'd236;
    mem[2385] = 'd232;
    mem[2386] = 'd224;
    mem[2387] = 'd220;
    mem[2388] = 'd148;
    mem[2389] = 'd144;
    mem[2390] = 'd84;
    mem[2391] = 'd84;
    mem[2392] = 'd264;
    mem[2393] = 'd320;
    mem[2394] = 'd188;
    mem[2395] = 'd220;
    mem[2396] = 'd84;
    mem[2397] = 'd84;
    mem[2398] = 'd152;
    mem[2399] = 'd148;
    mem[2400] = 'd184;
    mem[2401] = 'd180;
    mem[2402] = 'd188;
    mem[2403] = 'd180;
    mem[2404] = 'd188;
    mem[2405] = 'd188;
    mem[2406] = 'd196;
    mem[2407] = 'd192;
    mem[2408] = 'd200;
    mem[2409] = 'd196;
    mem[2410] = 'd188;
    mem[2411] = 'd184;
    mem[2412] = 'd172;
    mem[2413] = 'd168;
    mem[2414] = 'd156;
    mem[2415] = 'd148;
    mem[2416] = 'd140;
    mem[2417] = 'd140;
    mem[2418] = 'd104;
    mem[2419] = 'd104;
    mem[2420] = 'd88;
    mem[2421] = 'd88;
    mem[2422] = 'd420;
    mem[2423] = 'd600;
    mem[2424] = 'd612;
    mem[2425] = 'd908;
    mem[2426] = 'd572;
    mem[2427] = 'd948;
    mem[2428] = 'd692;
    mem[2429] = 'd940;
    mem[2430] = 'd1020;
    mem[2431] = 'd1020;
    mem[2432] = 'd1020;
    mem[2433] = 'd1020;
    mem[2434] = 'd288;
    mem[2435] = 'd616;
    mem[2436] = 'd24;
    mem[2437] = 'd588;
    mem[2438] = 'd76;
    mem[2439] = 'd652;
    mem[2440] = 'd84;
    mem[2441] = 'd540;
    mem[2442] = 'd92;
    mem[2443] = 'd96;
    mem[2444] = 'd88;
    mem[2445] = 'd88;
    mem[2446] = 'd104;
    mem[2447] = 'd104;
    mem[2448] = 'd112;
    mem[2449] = 'd116;
    mem[2450] = 'd124;
    mem[2451] = 'd128;
    mem[2452] = 'd136;
    mem[2453] = 'd144;
    mem[2454] = 'd148;
    mem[2455] = 'd156;
    mem[2456] = 'd148;
    mem[2457] = 'd152;
    mem[2458] = 'd144;
    mem[2459] = 'd148;
    mem[2460] = 'd148;
    mem[2461] = 'd152;
    mem[2462] = 'd128;
    mem[2463] = 'd132;
    mem[2464] = 'd108;
    mem[2465] = 'd108;
    mem[2466] = 'd80;
    mem[2467] = 'd80;
    mem[2468] = 'd136;
    mem[2469] = 'd704;
    mem[2470] = 'd124;
    mem[2471] = 'd568;
    mem[2472] = 'd84;
    mem[2473] = 'd84;
    mem[2474] = 'd116;
    mem[2475] = 'd120;
    mem[2476] = 'd160;
    mem[2477] = 'd168;
    mem[2478] = 'd176;
    mem[2479] = 'd180;
    mem[2480] = 'd180;
    mem[2481] = 'd184;
    mem[2482] = 'd192;
    mem[2483] = 'd196;
    mem[2484] = 'd196;
    mem[2485] = 'd204;
    mem[2486] = 'd188;
    mem[2487] = 'd196;
    mem[2488] = 'd180;
    mem[2489] = 'd184;
    mem[2490] = 'd172;
    mem[2491] = 'd176;
    mem[2492] = 'd160;
    mem[2493] = 'd160;
    mem[2494] = 'd124;
    mem[2495] = 'd128;
    mem[2496] = 'd96;
    mem[2497] = 'd108;
    mem[2498] = 'd44;
    mem[2499] = 'd552;
    mem[2500] = 'd68;
    mem[2501] = 'd636;
    mem[2502] = 'd28;
    mem[2503] = 'd588;
    mem[2504] = 'd240;
    mem[2505] = 'd600;
    mem[2506] = 'd1020;
    mem[2507] = 'd1020;
    mem[2508] = 'd1020;
    mem[2509] = 'd1020;
    mem[2510] = 'd616;
    mem[2511] = 'd920;
    mem[2512] = 'd588;
    mem[2513] = 'd956;
    mem[2514] = 'd652;
    mem[2515] = 'd960;
    mem[2516] = 'd540;
    mem[2517] = 'd768;
    mem[2518] = 'd96;
    mem[2519] = 'd96;
    mem[2520] = 'd88;
    mem[2521] = 'd88;
    mem[2522] = 'd104;
    mem[2523] = 'd104;
    mem[2524] = 'd116;
    mem[2525] = 'd112;
    mem[2526] = 'd128;
    mem[2527] = 'd124;
    mem[2528] = 'd144;
    mem[2529] = 'd140;
    mem[2530] = 'd156;
    mem[2531] = 'd148;
    mem[2532] = 'd152;
    mem[2533] = 'd148;
    mem[2534] = 'd148;
    mem[2535] = 'd144;
    mem[2536] = 'd152;
    mem[2537] = 'd148;
    mem[2538] = 'd132;
    mem[2539] = 'd128;
    mem[2540] = 'd108;
    mem[2541] = 'd108;
    mem[2542] = 'd80;
    mem[2543] = 'd76;
    mem[2544] = 'd704;
    mem[2545] = 'd844;
    mem[2546] = 'd568;
    mem[2547] = 'd672;
    mem[2548] = 'd84;
    mem[2549] = 'd80;
    mem[2550] = 'd120;
    mem[2551] = 'd120;
    mem[2552] = 'd168;
    mem[2553] = 'd164;
    mem[2554] = 'd180;
    mem[2555] = 'd172;
    mem[2556] = 'd184;
    mem[2557] = 'd180;
    mem[2558] = 'd196;
    mem[2559] = 'd192;
    mem[2560] = 'd204;
    mem[2561] = 'd200;
    mem[2562] = 'd196;
    mem[2563] = 'd192;
    mem[2564] = 'd184;
    mem[2565] = 'd180;
    mem[2566] = 'd176;
    mem[2567] = 'd172;
    mem[2568] = 'd160;
    mem[2569] = 'd160;
    mem[2570] = 'd128;
    mem[2571] = 'd124;
    mem[2572] = 'd108;
    mem[2573] = 'd112;
    mem[2574] = 'd552;
    mem[2575] = 'd812;
    mem[2576] = 'd636;
    mem[2577] = 'd936;
    mem[2578] = 'd588;
    mem[2579] = 'd960;
    mem[2580] = 'd600;
    mem[2581] = 'd912;
    mem[2582] = 'd1020;
    mem[2583] = 'd1020;
    mem[2584] = 'd1020;
    mem[2585] = 'd1020;
    mem[2586] = 'd168;
    mem[2587] = 'd556;
    mem[2588] = 'd28;
    mem[2589] = 'd588;
    mem[2590] = 'd68;
    mem[2591] = 'd660;
    mem[2592] = 'd68;
    mem[2593] = 'd624;
    mem[2594] = 'd88;
    mem[2595] = 'd192;
    mem[2596] = 'd108;
    mem[2597] = 'd108;
    mem[2598] = 'd132;
    mem[2599] = 'd136;
    mem[2600] = 'd164;
    mem[2601] = 'd168;
    mem[2602] = 'd176;
    mem[2603] = 'd180;
    mem[2604] = 'd180;
    mem[2605] = 'd184;
    mem[2606] = 'd180;
    mem[2607] = 'd184;
    mem[2608] = 'd184;
    mem[2609] = 'd192;
    mem[2610] = 'd188;
    mem[2611] = 'd196;
    mem[2612] = 'd180;
    mem[2613] = 'd184;
    mem[2614] = 'd128;
    mem[2615] = 'd132;
    mem[2616] = 'd116;
    mem[2617] = 'd120;
    mem[2618] = 'd88;
    mem[2619] = 'd260;
    mem[2620] = 'd180;
    mem[2621] = 'd876;
    mem[2622] = 'd168;
    mem[2623] = 'd848;
    mem[2624] = 'd80;
    mem[2625] = 'd156;
    mem[2626] = 'd120;
    mem[2627] = 'd120;
    mem[2628] = 'd172;
    mem[2629] = 'd176;
    mem[2630] = 'd208;
    mem[2631] = 'd212;
    mem[2632] = 'd212;
    mem[2633] = 'd216;
    mem[2634] = 'd208;
    mem[2635] = 'd212;
    mem[2636] = 'd204;
    mem[2637] = 'd212;
    mem[2638] = 'd212;
    mem[2639] = 'd216;
    mem[2640] = 'd212;
    mem[2641] = 'd216;
    mem[2642] = 'd200;
    mem[2643] = 'd204;
    mem[2644] = 'd160;
    mem[2645] = 'd164;
    mem[2646] = 'd136;
    mem[2647] = 'd136;
    mem[2648] = 'd76;
    mem[2649] = 'd224;
    mem[2650] = 'd40;
    mem[2651] = 'd596;
    mem[2652] = 'd68;
    mem[2653] = 'd652;
    mem[2654] = 'd32;
    mem[2655] = 'd592;
    mem[2656] = 'd136;
    mem[2657] = 'd540;
    mem[2658] = 'd1020;
    mem[2659] = 'd1020;
    mem[2660] = 'd1020;
    mem[2661] = 'd1020;
    mem[2662] = 'd556;
    mem[2663] = 'd896;
    mem[2664] = 'd588;
    mem[2665] = 'd956;
    mem[2666] = 'd660;
    mem[2667] = 'd972;
    mem[2668] = 'd624;
    mem[2669] = 'd904;
    mem[2670] = 'd192;
    mem[2671] = 'd240;
    mem[2672] = 'd108;
    mem[2673] = 'd108;
    mem[2674] = 'd136;
    mem[2675] = 'd132;
    mem[2676] = 'd168;
    mem[2677] = 'd164;
    mem[2678] = 'd180;
    mem[2679] = 'd176;
    mem[2680] = 'd184;
    mem[2681] = 'd180;
    mem[2682] = 'd184;
    mem[2683] = 'd180;
    mem[2684] = 'd192;
    mem[2685] = 'd188;
    mem[2686] = 'd196;
    mem[2687] = 'd192;
    mem[2688] = 'd184;
    mem[2689] = 'd180;
    mem[2690] = 'd132;
    mem[2691] = 'd128;
    mem[2692] = 'd120;
    mem[2693] = 'd116;
    mem[2694] = 'd260;
    mem[2695] = 'd296;
    mem[2696] = 'd876;
    mem[2697] = 'd1004;
    mem[2698] = 'd848;
    mem[2699] = 'd980;
    mem[2700] = 'd156;
    mem[2701] = 'd176;
    mem[2702] = 'd120;
    mem[2703] = 'd120;
    mem[2704] = 'd176;
    mem[2705] = 'd172;
    mem[2706] = 'd212;
    mem[2707] = 'd208;
    mem[2708] = 'd216;
    mem[2709] = 'd212;
    mem[2710] = 'd212;
    mem[2711] = 'd208;
    mem[2712] = 'd212;
    mem[2713] = 'd204;
    mem[2714] = 'd216;
    mem[2715] = 'd212;
    mem[2716] = 'd216;
    mem[2717] = 'd216;
    mem[2718] = 'd204;
    mem[2719] = 'd200;
    mem[2720] = 'd164;
    mem[2721] = 'd160;
    mem[2722] = 'd136;
    mem[2723] = 'd136;
    mem[2724] = 'd224;
    mem[2725] = 'd304;
    mem[2726] = 'd596;
    mem[2727] = 'd880;
    mem[2728] = 'd652;
    mem[2729] = 'd960;
    mem[2730] = 'd592;
    mem[2731] = 'd956;
    mem[2732] = 'd540;
    mem[2733] = 'd892;
    mem[2734] = 'd1020;
    mem[2735] = 'd1020;
    mem[2736] = 'd1020;
    mem[2737] = 'd1020;
    mem[2738] = 'd124;
    mem[2739] = 'd528;
    mem[2740] = 'd28;
    mem[2741] = 'd584;
    mem[2742] = 'd60;
    mem[2743] = 'd664;
    mem[2744] = 'd72;
    mem[2745] = 'd648;
    mem[2746] = 'd76;
    mem[2747] = 'd408;
    mem[2748] = 'd120;
    mem[2749] = 'd120;
    mem[2750] = 'd120;
    mem[2751] = 'd124;
    mem[2752] = 'd168;
    mem[2753] = 'd168;
    mem[2754] = 'd188;
    mem[2755] = 'd188;
    mem[2756] = 'd192;
    mem[2757] = 'd192;
    mem[2758] = 'd192;
    mem[2759] = 'd196;
    mem[2760] = 'd192;
    mem[2761] = 'd200;
    mem[2762] = 'd188;
    mem[2763] = 'd188;
    mem[2764] = 'd140;
    mem[2765] = 'd144;
    mem[2766] = 'd124;
    mem[2767] = 'd124;
    mem[2768] = 'd88;
    mem[2769] = 'd84;
    mem[2770] = 'd136;
    mem[2771] = 'd644;
    mem[2772] = 'd192;
    mem[2773] = 'd888;
    mem[2774] = 'd188;
    mem[2775] = 'd880;
    mem[2776] = 'd120;
    mem[2777] = 'd540;
    mem[2778] = 'd100;
    mem[2779] = 'd96;
    mem[2780] = 'd128;
    mem[2781] = 'd132;
    mem[2782] = 'd176;
    mem[2783] = 'd180;
    mem[2784] = 'd204;
    mem[2785] = 'd208;
    mem[2786] = 'd204;
    mem[2787] = 'd208;
    mem[2788] = 'd200;
    mem[2789] = 'd208;
    mem[2790] = 'd204;
    mem[2791] = 'd208;
    mem[2792] = 'd204;
    mem[2793] = 'd208;
    mem[2794] = 'd176;
    mem[2795] = 'd180;
    mem[2796] = 'd116;
    mem[2797] = 'd120;
    mem[2798] = 'd120;
    mem[2799] = 'd116;
    mem[2800] = 'd48;
    mem[2801] = 'd444;
    mem[2802] = 'd56;
    mem[2803] = 'd620;
    mem[2804] = 'd64;
    mem[2805] = 'd664;
    mem[2806] = 'd28;
    mem[2807] = 'd588;
    mem[2808] = 'd88;
    mem[2809] = 'd512;
    mem[2810] = 'd1012;
    mem[2811] = 'd1012;
    mem[2812] = 'd1020;
    mem[2813] = 'd1020;
    mem[2814] = 'd528;
    mem[2815] = 'd880;
    mem[2816] = 'd584;
    mem[2817] = 'd948;
    mem[2818] = 'd664;
    mem[2819] = 'd980;
    mem[2820] = 'd648;
    mem[2821] = 'd940;
    mem[2822] = 'd408;
    mem[2823] = 'd572;
    mem[2824] = 'd120;
    mem[2825] = 'd120;
    mem[2826] = 'd124;
    mem[2827] = 'd120;
    mem[2828] = 'd168;
    mem[2829] = 'd168;
    mem[2830] = 'd188;
    mem[2831] = 'd188;
    mem[2832] = 'd192;
    mem[2833] = 'd192;
    mem[2834] = 'd196;
    mem[2835] = 'd192;
    mem[2836] = 'd200;
    mem[2837] = 'd196;
    mem[2838] = 'd188;
    mem[2839] = 'd188;
    mem[2840] = 'd144;
    mem[2841] = 'd140;
    mem[2842] = 'd124;
    mem[2843] = 'd124;
    mem[2844] = 'd84;
    mem[2845] = 'd84;
    mem[2846] = 'd644;
    mem[2847] = 'd752;
    mem[2848] = 'd888;
    mem[2849] = 'd1016;
    mem[2850] = 'd880;
    mem[2851] = 'd1012;
    mem[2852] = 'd540;
    mem[2853] = 'd636;
    mem[2854] = 'd96;
    mem[2855] = 'd96;
    mem[2856] = 'd132;
    mem[2857] = 'd128;
    mem[2858] = 'd180;
    mem[2859] = 'd176;
    mem[2860] = 'd208;
    mem[2861] = 'd204;
    mem[2862] = 'd208;
    mem[2863] = 'd208;
    mem[2864] = 'd208;
    mem[2865] = 'd204;
    mem[2866] = 'd208;
    mem[2867] = 'd208;
    mem[2868] = 'd208;
    mem[2869] = 'd204;
    mem[2870] = 'd180;
    mem[2871] = 'd176;
    mem[2872] = 'd120;
    mem[2873] = 'd116;
    mem[2874] = 'd116;
    mem[2875] = 'd112;
    mem[2876] = 'd444;
    mem[2877] = 'd648;
    mem[2878] = 'd620;
    mem[2879] = 'd904;
    mem[2880] = 'd664;
    mem[2881] = 'd980;
    mem[2882] = 'd588;
    mem[2883] = 'd948;
    mem[2884] = 'd512;
    mem[2885] = 'd876;
    mem[2886] = 'd1012;
    mem[2887] = 'd1016;
    mem[2888] = 'd1020;
    mem[2889] = 'd1020;
    mem[2890] = 'd120;
    mem[2891] = 'd520;
    mem[2892] = 'd28;
    mem[2893] = 'd576;
    mem[2894] = 'd56;
    mem[2895] = 'd660;
    mem[2896] = 'd92;
    mem[2897] = 'd684;
    mem[2898] = 'd72;
    mem[2899] = 'd608;
    mem[2900] = 'd92;
    mem[2901] = 'd200;
    mem[2902] = 'd128;
    mem[2903] = 'd132;
    mem[2904] = 'd108;
    mem[2905] = 'd112;
    mem[2906] = 'd120;
    mem[2907] = 'd124;
    mem[2908] = 'd136;
    mem[2909] = 'd140;
    mem[2910] = 'd144;
    mem[2911] = 'd148;
    mem[2912] = 'd140;
    mem[2913] = 'd140;
    mem[2914] = 'd112;
    mem[2915] = 'd116;
    mem[2916] = 'd112;
    mem[2917] = 'd116;
    mem[2918] = 'd104;
    mem[2919] = 'd104;
    mem[2920] = 'd92;
    mem[2921] = 'd356;
    mem[2922] = 'd176;
    mem[2923] = 'd856;
    mem[2924] = 'd196;
    mem[2925] = 'd884;
    mem[2926] = 'd192;
    mem[2927] = 'd884;
    mem[2928] = 'd172;
    mem[2929] = 'd840;
    mem[2930] = 'd80;
    mem[2931] = 'd268;
    mem[2932] = 'd120;
    mem[2933] = 'd120;
    mem[2934] = 'd120;
    mem[2935] = 'd120;
    mem[2936] = 'd120;
    mem[2937] = 'd124;
    mem[2938] = 'd128;
    mem[2939] = 'd132;
    mem[2940] = 'd132;
    mem[2941] = 'd136;
    mem[2942] = 'd136;
    mem[2943] = 'd136;
    mem[2944] = 'd124;
    mem[2945] = 'd128;
    mem[2946] = 'd100;
    mem[2947] = 'd100;
    mem[2948] = 'd124;
    mem[2949] = 'd128;
    mem[2950] = 'd68;
    mem[2951] = 'd220;
    mem[2952] = 'd40;
    mem[2953] = 'd588;
    mem[2954] = 'd84;
    mem[2955] = 'd668;
    mem[2956] = 'd60;
    mem[2957] = 'd668;
    mem[2958] = 'd28;
    mem[2959] = 'd580;
    mem[2960] = 'd88;
    mem[2961] = 'd504;
    mem[2962] = 'd1012;
    mem[2963] = 'd1012;
    mem[2964] = 'd1020;
    mem[2965] = 'd1020;
    mem[2966] = 'd520;
    mem[2967] = 'd872;
    mem[2968] = 'd576;
    mem[2969] = 'd932;
    mem[2970] = 'd660;
    mem[2971] = 'd984;
    mem[2972] = 'd684;
    mem[2973] = 'd968;
    mem[2974] = 'd608;
    mem[2975] = 'd876;
    mem[2976] = 'd200;
    mem[2977] = 'd256;
    mem[2978] = 'd132;
    mem[2979] = 'd128;
    mem[2980] = 'd112;
    mem[2981] = 'd112;
    mem[2982] = 'd124;
    mem[2983] = 'd120;
    mem[2984] = 'd140;
    mem[2985] = 'd140;
    mem[2986] = 'd148;
    mem[2987] = 'd144;
    mem[2988] = 'd140;
    mem[2989] = 'd140;
    mem[2990] = 'd116;
    mem[2991] = 'd112;
    mem[2992] = 'd116;
    mem[2993] = 'd112;
    mem[2994] = 'd104;
    mem[2995] = 'd100;
    mem[2996] = 'd356;
    mem[2997] = 'd432;
    mem[2998] = 'd856;
    mem[2999] = 'd1008;
    mem[3000] = 'd884;
    mem[3001] = 'd1020;
    mem[3002] = 'd884;
    mem[3003] = 'd1020;
    mem[3004] = 'd840;
    mem[3005] = 'd992;
    mem[3006] = 'd268;
    mem[3007] = 'd324;
    mem[3008] = 'd120;
    mem[3009] = 'd120;
    mem[3010] = 'd120;
    mem[3011] = 'd120;
    mem[3012] = 'd124;
    mem[3013] = 'd120;
    mem[3014] = 'd132;
    mem[3015] = 'd132;
    mem[3016] = 'd136;
    mem[3017] = 'd136;
    mem[3018] = 'd136;
    mem[3019] = 'd132;
    mem[3020] = 'd128;
    mem[3021] = 'd124;
    mem[3022] = 'd100;
    mem[3023] = 'd100;
    mem[3024] = 'd128;
    mem[3025] = 'd128;
    mem[3026] = 'd220;
    mem[3027] = 'd300;
    mem[3028] = 'd588;
    mem[3029] = 'd872;
    mem[3030] = 'd668;
    mem[3031] = 'd956;
    mem[3032] = 'd668;
    mem[3033] = 'd984;
    mem[3034] = 'd580;
    mem[3035] = 'd940;
    mem[3036] = 'd504;
    mem[3037] = 'd872;
    mem[3038] = 'd1012;
    mem[3039] = 'd1016;
    mem[3040] = 'd1020;
    mem[3041] = 'd1020;
    mem[3042] = 'd168;
    mem[3043] = 'd536;
    mem[3044] = 'd24;
    mem[3045] = 'd560;
    mem[3046] = 'd48;
    mem[3047] = 'd648;
    mem[3048] = 'd104;
    mem[3049] = 'd700;
    mem[3050] = 'd112;
    mem[3051] = 'd680;
    mem[3052] = 'd76;
    mem[3053] = 'd548;
    mem[3054] = 'd84;
    mem[3055] = 'd168;
    mem[3056] = 'd132;
    mem[3057] = 'd132;
    mem[3058] = 'd152;
    mem[3059] = 'd152;
    mem[3060] = 'd152;
    mem[3061] = 'd152;
    mem[3062] = 'd152;
    mem[3063] = 'd156;
    mem[3064] = 'd144;
    mem[3065] = 'd144;
    mem[3066] = 'd136;
    mem[3067] = 'd136;
    mem[3068] = 'd88;
    mem[3069] = 'd88;
    mem[3070] = 'd84;
    mem[3071] = 'd360;
    mem[3072] = 'd164;
    mem[3073] = 'd816;
    mem[3074] = 'd196;
    mem[3075] = 'd868;
    mem[3076] = 'd200;
    mem[3077] = 'd876;
    mem[3078] = 'd196;
    mem[3079] = 'd876;
    mem[3080] = 'd196;
    mem[3081] = 'd868;
    mem[3082] = 'd152;
    mem[3083] = 'd780;
    mem[3084] = 'd76;
    mem[3085] = 'd288;
    mem[3086] = 'd104;
    mem[3087] = 'd100;
    mem[3088] = 'd156;
    mem[3089] = 'd156;
    mem[3090] = 'd152;
    mem[3091] = 'd152;
    mem[3092] = 'd148;
    mem[3093] = 'd152;
    mem[3094] = 'd144;
    mem[3095] = 'd148;
    mem[3096] = 'd140;
    mem[3097] = 'd144;
    mem[3098] = 'd132;
    mem[3099] = 'd128;
    mem[3100] = 'd68;
    mem[3101] = 'd164;
    mem[3102] = 'd44;
    mem[3103] = 'd556;
    mem[3104] = 'd96;
    mem[3105] = 'd660;
    mem[3106] = 'd100;
    mem[3107] = 'd700;
    mem[3108] = 'd52;
    mem[3109] = 'd652;
    mem[3110] = 'd28;
    mem[3111] = 'd568;
    mem[3112] = 'd136;
    mem[3113] = 'd520;
    mem[3114] = 'd1020;
    mem[3115] = 'd1020;
    mem[3116] = 'd1020;
    mem[3117] = 'd1020;
    mem[3118] = 'd536;
    mem[3119] = 'd868;
    mem[3120] = 'd560;
    mem[3121] = 'd924;
    mem[3122] = 'd648;
    mem[3123] = 'd976;
    mem[3124] = 'd700;
    mem[3125] = 'd996;
    mem[3126] = 'd680;
    mem[3127] = 'd956;
    mem[3128] = 'd548;
    mem[3129] = 'd780;
    mem[3130] = 'd168;
    mem[3131] = 'd208;
    mem[3132] = 'd132;
    mem[3133] = 'd128;
    mem[3134] = 'd152;
    mem[3135] = 'd152;
    mem[3136] = 'd152;
    mem[3137] = 'd152;
    mem[3138] = 'd156;
    mem[3139] = 'd152;
    mem[3140] = 'd144;
    mem[3141] = 'd144;
    mem[3142] = 'd136;
    mem[3143] = 'd136;
    mem[3144] = 'd88;
    mem[3145] = 'd88;
    mem[3146] = 'd360;
    mem[3147] = 'd452;
    mem[3148] = 'd816;
    mem[3149] = 'd984;
    mem[3150] = 'd868;
    mem[3151] = 'd1016;
    mem[3152] = 'd876;
    mem[3153] = 'd1020;
    mem[3154] = 'd876;
    mem[3155] = 'd1020;
    mem[3156] = 'd868;
    mem[3157] = 'd1016;
    mem[3158] = 'd780;
    mem[3159] = 'd956;
    mem[3160] = 'd288;
    mem[3161] = 'd356;
    mem[3162] = 'd100;
    mem[3163] = 'd100;
    mem[3164] = 'd156;
    mem[3165] = 'd156;
    mem[3166] = 'd152;
    mem[3167] = 'd152;
    mem[3168] = 'd152;
    mem[3169] = 'd148;
    mem[3170] = 'd148;
    mem[3171] = 'd144;
    mem[3172] = 'd144;
    mem[3173] = 'd140;
    mem[3174] = 'd128;
    mem[3175] = 'd124;
    mem[3176] = 'd164;
    mem[3177] = 'd216;
    mem[3178] = 'd556;
    mem[3179] = 'd816;
    mem[3180] = 'd660;
    mem[3181] = 'd936;
    mem[3182] = 'd700;
    mem[3183] = 'd996;
    mem[3184] = 'd652;
    mem[3185] = 'd980;
    mem[3186] = 'd568;
    mem[3187] = 'd928;
    mem[3188] = 'd520;
    mem[3189] = 'd864;
    mem[3190] = 'd1020;
    mem[3191] = 'd1020;
    mem[3192] = 'd1020;
    mem[3193] = 'd1020;
    mem[3194] = 'd280;
    mem[3195] = 'd592;
    mem[3196] = 'd24;
    mem[3197] = 'd540;
    mem[3198] = 'd44;
    mem[3199] = 'd632;
    mem[3200] = 'd88;
    mem[3201] = 'd700;
    mem[3202] = 'd140;
    mem[3203] = 'd728;
    mem[3204] = 'd144;
    mem[3205] = 'd708;
    mem[3206] = 'd108;
    mem[3207] = 'd640;
    mem[3208] = 'd84;
    mem[3209] = 'd440;
    mem[3210] = 'd76;
    mem[3211] = 'd268;
    mem[3212] = 'd72;
    mem[3213] = 'd184;
    mem[3214] = 'd72;
    mem[3215] = 'd156;
    mem[3216] = 'd72;
    mem[3217] = 'd204;
    mem[3218] = 'd88;
    mem[3219] = 'd336;
    mem[3220] = 'd132;
    mem[3221] = 'd636;
    mem[3222] = 'd184;
    mem[3223] = 'd828;
    mem[3224] = 'd208;
    mem[3225] = 'd856;
    mem[3226] = 'd208;
    mem[3227] = 'd864;
    mem[3228] = 'd204;
    mem[3229] = 'd864;
    mem[3230] = 'd208;
    mem[3231] = 'd864;
    mem[3232] = 'd208;
    mem[3233] = 'd864;
    mem[3234] = 'd204;
    mem[3235] = 'd856;
    mem[3236] = 'd176;
    mem[3237] = 'd812;
    mem[3238] = 'd108;
    mem[3239] = 'd572;
    mem[3240] = 'd72;
    mem[3241] = 'd292;
    mem[3242] = 'd64;
    mem[3243] = 'd188;
    mem[3244] = 'd64;
    mem[3245] = 'd148;
    mem[3246] = 'd64;
    mem[3247] = 'd176;
    mem[3248] = 'd60;
    mem[3249] = 'd276;
    mem[3250] = 'd60;
    mem[3251] = 'd428;
    mem[3252] = 'd76;
    mem[3253] = 'd632;
    mem[3254] = 'd132;
    mem[3255] = 'd692;
    mem[3256] = 'd140;
    mem[3257] = 'd724;
    mem[3258] = 'd84;
    mem[3259] = 'd700;
    mem[3260] = 'd48;
    mem[3261] = 'd636;
    mem[3262] = 'd28;
    mem[3263] = 'd548;
    mem[3264] = 'd236;
    mem[3265] = 'd568;
    mem[3266] = 'd1020;
    mem[3267] = 'd1020;
    mem[3268] = 'd1020;
    mem[3269] = 'd1020;
    mem[3270] = 'd592;
    mem[3271] = 'd876;
    mem[3272] = 'd540;
    mem[3273] = 'd908;
    mem[3274] = 'd632;
    mem[3275] = 'd960;
    mem[3276] = 'd700;
    mem[3277] = 'd1000;
    mem[3278] = 'd728;
    mem[3279] = 'd1004;
    mem[3280] = 'd708;
    mem[3281] = 'd976;
    mem[3282] = 'd640;
    mem[3283] = 'd888;
    mem[3284] = 'd440;
    mem[3285] = 'd604;
    mem[3286] = 'd268;
    mem[3287] = 'd360;
    mem[3288] = 'd184;
    mem[3289] = 'd228;
    mem[3290] = 'd156;
    mem[3291] = 'd192;
    mem[3292] = 'd204;
    mem[3293] = 'd260;
    mem[3294] = 'd336;
    mem[3295] = 'd432;
    mem[3296] = 'd636;
    mem[3297] = 'd804;
    mem[3298] = 'd828;
    mem[3299] = 'd1004;
    mem[3300] = 'd856;
    mem[3301] = 'd1020;
    mem[3302] = 'd864;
    mem[3303] = 'd1020;
    mem[3304] = 'd864;
    mem[3305] = 'd1020;
    mem[3306] = 'd864;
    mem[3307] = 'd1020;
    mem[3308] = 'd864;
    mem[3309] = 'd1020;
    mem[3310] = 'd856;
    mem[3311] = 'd1016;
    mem[3312] = 'd812;
    mem[3313] = 'd996;
    mem[3314] = 'd572;
    mem[3315] = 'd736;
    mem[3316] = 'd292;
    mem[3317] = 'd376;
    mem[3318] = 'd188;
    mem[3319] = 'd244;
    mem[3320] = 'd148;
    mem[3321] = 'd188;
    mem[3322] = 'd176;
    mem[3323] = 'd232;
    mem[3324] = 'd276;
    mem[3325] = 'd384;
    mem[3326] = 'd428;
    mem[3327] = 'd604;
    mem[3328] = 'd632;
    mem[3329] = 'd900;
    mem[3330] = 'd692;
    mem[3331] = 'd956;
    mem[3332] = 'd724;
    mem[3333] = 'd1004;
    mem[3334] = 'd700;
    mem[3335] = 'd1004;
    mem[3336] = 'd636;
    mem[3337] = 'd964;
    mem[3338] = 'd548;
    mem[3339] = 'd912;
    mem[3340] = 'd568;
    mem[3341] = 'd872;
    mem[3342] = 'd1020;
    mem[3343] = 'd1020;
    mem[3344] = 'd1020;
    mem[3345] = 'd1020;
    mem[3346] = 'd448;
    mem[3347] = 'd676;
    mem[3348] = 'd20;
    mem[3349] = 'd516;
    mem[3350] = 'd44;
    mem[3351] = 'd612;
    mem[3352] = 'd68;
    mem[3353] = 'd684;
    mem[3354] = 'd120;
    mem[3355] = 'd720;
    mem[3356] = 'd172;
    mem[3357] = 'd744;
    mem[3358] = 'd188;
    mem[3359] = 'd760;
    mem[3360] = 'd180;
    mem[3361] = 'd760;
    mem[3362] = 'd172;
    mem[3363] = 'd756;
    mem[3364] = 'd160;
    mem[3365] = 'd756;
    mem[3366] = 'd164;
    mem[3367] = 'd768;
    mem[3368] = 'd176;
    mem[3369] = 'd788;
    mem[3370] = 'd196;
    mem[3371] = 'd812;
    mem[3372] = 'd204;
    mem[3373] = 'd836;
    mem[3374] = 'd208;
    mem[3375] = 'd844;
    mem[3376] = 'd212;
    mem[3377] = 'd848;
    mem[3378] = 'd208;
    mem[3379] = 'd852;
    mem[3380] = 'd208;
    mem[3381] = 'd852;
    mem[3382] = 'd208;
    mem[3383] = 'd852;
    mem[3384] = 'd208;
    mem[3385] = 'd852;
    mem[3386] = 'd208;
    mem[3387] = 'd852;
    mem[3388] = 'd208;
    mem[3389] = 'd844;
    mem[3390] = 'd200;
    mem[3391] = 'd832;
    mem[3392] = 'd184;
    mem[3393] = 'd800;
    mem[3394] = 'd160;
    mem[3395] = 'd764;
    mem[3396] = 'd148;
    mem[3397] = 'd744;
    mem[3398] = 'd148;
    mem[3399] = 'd736;
    mem[3400] = 'd160;
    mem[3401] = 'd740;
    mem[3402] = 'd172;
    mem[3403] = 'd748;
    mem[3404] = 'd188;
    mem[3405] = 'd756;
    mem[3406] = 'd172;
    mem[3407] = 'd748;
    mem[3408] = 'd120;
    mem[3409] = 'd724;
    mem[3410] = 'd72;
    mem[3411] = 'd684;
    mem[3412] = 'd48;
    mem[3413] = 'd616;
    mem[3414] = 'd24;
    mem[3415] = 'd524;
    mem[3416] = 'd404;
    mem[3417] = 'd660;
    mem[3418] = 'd1020;
    mem[3419] = 'd1020;
    mem[3420] = 'd1020;
    mem[3421] = 'd1020;
    mem[3422] = 'd676;
    mem[3423] = 'd900;
    mem[3424] = 'd516;
    mem[3425] = 'd884;
    mem[3426] = 'd612;
    mem[3427] = 'd944;
    mem[3428] = 'd684;
    mem[3429] = 'd996;
    mem[3430] = 'd720;
    mem[3431] = 'd1012;
    mem[3432] = 'd744;
    mem[3433] = 'd1016;
    mem[3434] = 'd760;
    mem[3435] = 'd1012;
    mem[3436] = 'd760;
    mem[3437] = 'd1000;
    mem[3438] = 'd756;
    mem[3439] = 'd988;
    mem[3440] = 'd756;
    mem[3441] = 'd988;
    mem[3442] = 'd768;
    mem[3443] = 'd992;
    mem[3444] = 'd788;
    mem[3445] = 'd1000;
    mem[3446] = 'd812;
    mem[3447] = 'd1008;
    mem[3448] = 'd836;
    mem[3449] = 'd1016;
    mem[3450] = 'd844;
    mem[3451] = 'd1020;
    mem[3452] = 'd848;
    mem[3453] = 'd1020;
    mem[3454] = 'd852;
    mem[3455] = 'd1020;
    mem[3456] = 'd852;
    mem[3457] = 'd1020;
    mem[3458] = 'd852;
    mem[3459] = 'd1020;
    mem[3460] = 'd852;
    mem[3461] = 'd1020;
    mem[3462] = 'd852;
    mem[3463] = 'd1020;
    mem[3464] = 'd844;
    mem[3465] = 'd1020;
    mem[3466] = 'd832;
    mem[3467] = 'd1012;
    mem[3468] = 'd800;
    mem[3469] = 'd996;
    mem[3470] = 'd764;
    mem[3471] = 'd984;
    mem[3472] = 'd744;
    mem[3473] = 'd976;
    mem[3474] = 'd736;
    mem[3475] = 'd972;
    mem[3476] = 'd740;
    mem[3477] = 'd976;
    mem[3478] = 'd748;
    mem[3479] = 'd992;
    mem[3480] = 'd756;
    mem[3481] = 'd1008;
    mem[3482] = 'd748;
    mem[3483] = 'd1016;
    mem[3484] = 'd724;
    mem[3485] = 'd1012;
    mem[3486] = 'd684;
    mem[3487] = 'd996;
    mem[3488] = 'd616;
    mem[3489] = 'd948;
    mem[3490] = 'd524;
    mem[3491] = 'd892;
    mem[3492] = 'd660;
    mem[3493] = 'd892;
    mem[3494] = 'd1020;
    mem[3495] = 'd1020;
    mem[3496] = 'd1020;
    mem[3497] = 'd1020;
    mem[3498] = 'd676;
    mem[3499] = 'd808;
    mem[3500] = 'd16;
    mem[3501] = 'd488;
    mem[3502] = 'd40;
    mem[3503] = 'd584;
    mem[3504] = 'd64;
    mem[3505] = 'd660;
    mem[3506] = 'd92;
    mem[3507] = 'd704;
    mem[3508] = 'd140;
    mem[3509] = 'd732;
    mem[3510] = 'd184;
    mem[3511] = 'd756;
    mem[3512] = 'd208;
    mem[3513] = 'd772;
    mem[3514] = 'd212;
    mem[3515] = 'd784;
    mem[3516] = 'd200;
    mem[3517] = 'd780;
    mem[3518] = 'd204;
    mem[3519] = 'd800;
    mem[3520] = 'd212;
    mem[3521] = 'd816;
    mem[3522] = 'd216;
    mem[3523] = 'd824;
    mem[3524] = 'd216;
    mem[3525] = 'd832;
    mem[3526] = 'd216;
    mem[3527] = 'd836;
    mem[3528] = 'd216;
    mem[3529] = 'd836;
    mem[3530] = 'd216;
    mem[3531] = 'd840;
    mem[3532] = 'd220;
    mem[3533] = 'd840;
    mem[3534] = 'd216;
    mem[3535] = 'd844;
    mem[3536] = 'd216;
    mem[3537] = 'd840;
    mem[3538] = 'd216;
    mem[3539] = 'd836;
    mem[3540] = 'd216;
    mem[3541] = 'd836;
    mem[3542] = 'd216;
    mem[3543] = 'd832;
    mem[3544] = 'd216;
    mem[3545] = 'd824;
    mem[3546] = 'd216;
    mem[3547] = 'd820;
    mem[3548] = 'd208;
    mem[3549] = 'd800;
    mem[3550] = 'd200;
    mem[3551] = 'd776;
    mem[3552] = 'd212;
    mem[3553] = 'd784;
    mem[3554] = 'd208;
    mem[3555] = 'd772;
    mem[3556] = 'd184;
    mem[3557] = 'd756;
    mem[3558] = 'd144;
    mem[3559] = 'd732;
    mem[3560] = 'd92;
    mem[3561] = 'd708;
    mem[3562] = 'd64;
    mem[3563] = 'd660;
    mem[3564] = 'd44;
    mem[3565] = 'd588;
    mem[3566] = 'd16;
    mem[3567] = 'd492;
    mem[3568] = 'd636;
    mem[3569] = 'd788;
    mem[3570] = 'd1020;
    mem[3571] = 'd1020;
    mem[3572] = 'd1020;
    mem[3573] = 'd1020;
    mem[3574] = 'd808;
    mem[3575] = 'd936;
    mem[3576] = 'd488;
    mem[3577] = 'd860;
    mem[3578] = 'd584;
    mem[3579] = 'd924;
    mem[3580] = 'd660;
    mem[3581] = 'd976;
    mem[3582] = 'd704;
    mem[3583] = 'd1008;
    mem[3584] = 'd732;
    mem[3585] = 'd1016;
    mem[3586] = 'd756;
    mem[3587] = 'd1020;
    mem[3588] = 'd772;
    mem[3589] = 'd1020;
    mem[3590] = 'd784;
    mem[3591] = 'd1020;
    mem[3592] = 'd780;
    mem[3593] = 'd1008;
    mem[3594] = 'd800;
    mem[3595] = 'd1012;
    mem[3596] = 'd816;
    mem[3597] = 'd1020;
    mem[3598] = 'd824;
    mem[3599] = 'd1020;
    mem[3600] = 'd832;
    mem[3601] = 'd1020;
    mem[3602] = 'd836;
    mem[3603] = 'd1020;
    mem[3604] = 'd836;
    mem[3605] = 'd1020;
    mem[3606] = 'd840;
    mem[3607] = 'd1020;
    mem[3608] = 'd840;
    mem[3609] = 'd1020;
    mem[3610] = 'd844;
    mem[3611] = 'd1020;
    mem[3612] = 'd840;
    mem[3613] = 'd1020;
    mem[3614] = 'd836;
    mem[3615] = 'd1020;
    mem[3616] = 'd836;
    mem[3617] = 'd1020;
    mem[3618] = 'd832;
    mem[3619] = 'd1020;
    mem[3620] = 'd824;
    mem[3621] = 'd1020;
    mem[3622] = 'd820;
    mem[3623] = 'd1020;
    mem[3624] = 'd800;
    mem[3625] = 'd1016;
    mem[3626] = 'd776;
    mem[3627] = 'd1012;
    mem[3628] = 'd784;
    mem[3629] = 'd1020;
    mem[3630] = 'd772;
    mem[3631] = 'd1020;
    mem[3632] = 'd756;
    mem[3633] = 'd1020;
    mem[3634] = 'd732;
    mem[3635] = 'd1016;
    mem[3636] = 'd708;
    mem[3637] = 'd1008;
    mem[3638] = 'd660;
    mem[3639] = 'd976;
    mem[3640] = 'd588;
    mem[3641] = 'd928;
    mem[3642] = 'd492;
    mem[3643] = 'd864;
    mem[3644] = 'd788;
    mem[3645] = 'd928;
    mem[3646] = 'd1020;
    mem[3647] = 'd1020;
    mem[3648] = 'd1020;
    mem[3649] = 'd1020;
    mem[3650] = 'd944;
    mem[3651] = 'd968;
    mem[3652] = 'd36;
    mem[3653] = 'd460;
    mem[3654] = 'd36;
    mem[3655] = 'd548;
    mem[3656] = 'd56;
    mem[3657] = 'd636;
    mem[3658] = 'd76;
    mem[3659] = 'd684;
    mem[3660] = 'd108;
    mem[3661] = 'd716;
    mem[3662] = 'd156;
    mem[3663] = 'd740;
    mem[3664] = 'd196;
    mem[3665] = 'd756;
    mem[3666] = 'd216;
    mem[3667] = 'd772;
    mem[3668] = 'd112;
    mem[3669] = 'd480;
    mem[3670] = 'd104;
    mem[3671] = 'd500;
    mem[3672] = 'd200;
    mem[3673] = 'd776;
    mem[3674] = 'd216;
    mem[3675] = 'd812;
    mem[3676] = 'd224;
    mem[3677] = 'd820;
    mem[3678] = 'd220;
    mem[3679] = 'd824;
    mem[3680] = 'd224;
    mem[3681] = 'd828;
    mem[3682] = 'd220;
    mem[3683] = 'd828;
    mem[3684] = 'd220;
    mem[3685] = 'd828;
    mem[3686] = 'd220;
    mem[3687] = 'd828;
    mem[3688] = 'd220;
    mem[3689] = 'd828;
    mem[3690] = 'd220;
    mem[3691] = 'd828;
    mem[3692] = 'd220;
    mem[3693] = 'd824;
    mem[3694] = 'd220;
    mem[3695] = 'd820;
    mem[3696] = 'd220;
    mem[3697] = 'd812;
    mem[3698] = 'd200;
    mem[3699] = 'd772;
    mem[3700] = 'd84;
    mem[3701] = 'd436;
    mem[3702] = 'd136;
    mem[3703] = 'd544;
    mem[3704] = 'd216;
    mem[3705] = 'd772;
    mem[3706] = 'd196;
    mem[3707] = 'd756;
    mem[3708] = 'd156;
    mem[3709] = 'd736;
    mem[3710] = 'd112;
    mem[3711] = 'd720;
    mem[3712] = 'd76;
    mem[3713] = 'd684;
    mem[3714] = 'd60;
    mem[3715] = 'd636;
    mem[3716] = 'd36;
    mem[3717] = 'd556;
    mem[3718] = 'd24;
    mem[3719] = 'd464;
    mem[3720] = 'd916;
    mem[3721] = 'd952;
    mem[3722] = 'd1020;
    mem[3723] = 'd1020;
    mem[3724] = 'd1020;
    mem[3725] = 'd1020;
    mem[3726] = 'd968;
    mem[3727] = 'd996;
    mem[3728] = 'd460;
    mem[3729] = 'd832;
    mem[3730] = 'd548;
    mem[3731] = 'd896;
    mem[3732] = 'd636;
    mem[3733] = 'd956;
    mem[3734] = 'd684;
    mem[3735] = 'd996;
    mem[3736] = 'd716;
    mem[3737] = 'd1012;
    mem[3738] = 'd740;
    mem[3739] = 'd1016;
    mem[3740] = 'd756;
    mem[3741] = 'd1020;
    mem[3742] = 'd772;
    mem[3743] = 'd1020;
    mem[3744] = 'd480;
    mem[3745] = 'd704;
    mem[3746] = 'd500;
    mem[3747] = 'd748;
    mem[3748] = 'd776;
    mem[3749] = 'd1000;
    mem[3750] = 'd812;
    mem[3751] = 'd1020;
    mem[3752] = 'd820;
    mem[3753] = 'd1020;
    mem[3754] = 'd824;
    mem[3755] = 'd1020;
    mem[3756] = 'd828;
    mem[3757] = 'd1020;
    mem[3758] = 'd828;
    mem[3759] = 'd1020;
    mem[3760] = 'd828;
    mem[3761] = 'd1020;
    mem[3762] = 'd828;
    mem[3763] = 'd1020;
    mem[3764] = 'd828;
    mem[3765] = 'd1020;
    mem[3766] = 'd828;
    mem[3767] = 'd1020;
    mem[3768] = 'd824;
    mem[3769] = 'd1020;
    mem[3770] = 'd820;
    mem[3771] = 'd1020;
    mem[3772] = 'd812;
    mem[3773] = 'd1020;
    mem[3774] = 'd772;
    mem[3775] = 'd1000;
    mem[3776] = 'd436;
    mem[3777] = 'd680;
    mem[3778] = 'd544;
    mem[3779] = 'd760;
    mem[3780] = 'd772;
    mem[3781] = 'd1020;
    mem[3782] = 'd756;
    mem[3783] = 'd1020;
    mem[3784] = 'd736;
    mem[3785] = 'd1016;
    mem[3786] = 'd720;
    mem[3787] = 'd1012;
    mem[3788] = 'd684;
    mem[3789] = 'd1000;
    mem[3790] = 'd636;
    mem[3791] = 'd956;
    mem[3792] = 'd556;
    mem[3793] = 'd904;
    mem[3794] = 'd464;
    mem[3795] = 'd840;
    mem[3796] = 'd952;
    mem[3797] = 'd984;
    mem[3798] = 'd1020;
    mem[3799] = 'd1020;
    mem[3800] = 'd1020;
    mem[3801] = 'd1020;
    mem[3802] = 'd1020;
    mem[3803] = 'd1020;
    mem[3804] = 'd356;
    mem[3805] = 'd624;
    mem[3806] = 'd24;
    mem[3807] = 'd504;
    mem[3808] = 'd52;
    mem[3809] = 'd600;
    mem[3810] = 'd68;
    mem[3811] = 'd656;
    mem[3812] = 'd84;
    mem[3813] = 'd692;
    mem[3814] = 'd112;
    mem[3815] = 'd720;
    mem[3816] = 'd160;
    mem[3817] = 'd740;
    mem[3818] = 'd192;
    mem[3819] = 'd756;
    mem[3820] = 'd224;
    mem[3821] = 'd736;
    mem[3822] = 'd44;
    mem[3823] = 'd288;
    mem[3824] = 'd44;
    mem[3825] = 'd332;
    mem[3826] = 'd128;
    mem[3827] = 'd572;
    mem[3828] = 'd204;
    mem[3829] = 'd764;
    mem[3830] = 'd224;
    mem[3831] = 'd804;
    mem[3832] = 'd228;
    mem[3833] = 'd812;
    mem[3834] = 'd228;
    mem[3835] = 'd812;
    mem[3836] = 'd228;
    mem[3837] = 'd816;
    mem[3838] = 'd228;
    mem[3839] = 'd816;
    mem[3840] = 'd228;
    mem[3841] = 'd812;
    mem[3842] = 'd224;
    mem[3843] = 'd808;
    mem[3844] = 'd220;
    mem[3845] = 'd796;
    mem[3846] = 'd192;
    mem[3847] = 'd736;
    mem[3848] = 'd116;
    mem[3849] = 'd532;
    mem[3850] = 'd36;
    mem[3851] = 'd300;
    mem[3852] = 'd64;
    mem[3853] = 'd328;
    mem[3854] = 'd236;
    mem[3855] = 'd772;
    mem[3856] = 'd196;
    mem[3857] = 'd752;
    mem[3858] = 'd160;
    mem[3859] = 'd740;
    mem[3860] = 'd116;
    mem[3861] = 'd724;
    mem[3862] = 'd84;
    mem[3863] = 'd696;
    mem[3864] = 'd72;
    mem[3865] = 'd660;
    mem[3866] = 'd56;
    mem[3867] = 'd604;
    mem[3868] = 'd28;
    mem[3869] = 'd508;
    mem[3870] = 'd292;
    mem[3871] = 'd584;
    mem[3872] = 'd1020;
    mem[3873] = 'd1020;
    mem[3874] = 'd1020;
    mem[3875] = 'd1020;
    mem[3876] = 'd1020;
    mem[3877] = 'd1020;
    mem[3878] = 'd1020;
    mem[3879] = 'd1020;
    mem[3880] = 'd624;
    mem[3881] = 'd876;
    mem[3882] = 'd504;
    mem[3883] = 'd860;
    mem[3884] = 'd600;
    mem[3885] = 'd924;
    mem[3886] = 'd656;
    mem[3887] = 'd972;
    mem[3888] = 'd692;
    mem[3889] = 'd1004;
    mem[3890] = 'd720;
    mem[3891] = 'd1016;
    mem[3892] = 'd740;
    mem[3893] = 'd1016;
    mem[3894] = 'd756;
    mem[3895] = 'd1020;
    mem[3896] = 'd736;
    mem[3897] = 'd948;
    mem[3898] = 'd288;
    mem[3899] = 'd500;
    mem[3900] = 'd332;
    mem[3901] = 'd564;
    mem[3902] = 'd572;
    mem[3903] = 'd820;
    mem[3904] = 'd764;
    mem[3905] = 'd1000;
    mem[3906] = 'd804;
    mem[3907] = 'd1016;
    mem[3908] = 'd812;
    mem[3909] = 'd1020;
    mem[3910] = 'd812;
    mem[3911] = 'd1020;
    mem[3912] = 'd816;
    mem[3913] = 'd1020;
    mem[3914] = 'd816;
    mem[3915] = 'd1020;
    mem[3916] = 'd812;
    mem[3917] = 'd1020;
    mem[3918] = 'd808;
    mem[3919] = 'd1020;
    mem[3920] = 'd796;
    mem[3921] = 'd1016;
    mem[3922] = 'd736;
    mem[3923] = 'd972;
    mem[3924] = 'd532;
    mem[3925] = 'd780;
    mem[3926] = 'd300;
    mem[3927] = 'd528;
    mem[3928] = 'd328;
    mem[3929] = 'd528;
    mem[3930] = 'd772;
    mem[3931] = 'd988;
    mem[3932] = 'd752;
    mem[3933] = 'd1020;
    mem[3934] = 'd740;
    mem[3935] = 'd1016;
    mem[3936] = 'd724;
    mem[3937] = 'd1016;
    mem[3938] = 'd696;
    mem[3939] = 'd1004;
    mem[3940] = 'd660;
    mem[3941] = 'd972;
    mem[3942] = 'd604;
    mem[3943] = 'd928;
    mem[3944] = 'd508;
    mem[3945] = 'd868;
    mem[3946] = 'd584;
    mem[3947] = 'd864;
    mem[3948] = 'd1020;
    mem[3949] = 'd1020;
    mem[3950] = 'd1020;
    mem[3951] = 'd1020;
    mem[3952] = 'd1020;
    mem[3953] = 'd1020;
    mem[3954] = 'd1020;
    mem[3955] = 'd1020;
    mem[3956] = 'd792;
    mem[3957] = 'd876;
    mem[3958] = 'd12;
    mem[3959] = 'd456;
    mem[3960] = 'd40;
    mem[3961] = 'd556;
    mem[3962] = 'd64;
    mem[3963] = 'd624;
    mem[3964] = 'd80;
    mem[3965] = 'd668;
    mem[3966] = 'd88;
    mem[3967] = 'd700;
    mem[3968] = 'd116;
    mem[3969] = 'd716;
    mem[3970] = 'd156;
    mem[3971] = 'd736;
    mem[3972] = 'd192;
    mem[3973] = 'd752;
    mem[3974] = 'd216;
    mem[3975] = 'd712;
    mem[3976] = 'd48;
    mem[3977] = 'd332;
    mem[3978] = 'd20;
    mem[3979] = 'd252;
    mem[3980] = 'd32;
    mem[3981] = 'd288;
    mem[3982] = 'd76;
    mem[3983] = 'd420;
    mem[3984] = 'd120;
    mem[3985] = 'd548;
    mem[3986] = 'd152;
    mem[3987] = 'd640;
    mem[3988] = 'd168;
    mem[3989] = 'd676;
    mem[3990] = 'd164;
    mem[3991] = 'd672;
    mem[3992] = 'd152;
    mem[3993] = 'd628;
    mem[3994] = 'd116;
    mem[3995] = 'd536;
    mem[3996] = 'd72;
    mem[3997] = 'd404;
    mem[3998] = 'd32;
    mem[3999] = 'd288;
    mem[4000] = 'd16;
    mem[4001] = 'd256;
    mem[4002] = 'd68;
    mem[4003] = 'd372;
    mem[4004] = 'd232;
    mem[4005] = 'd752;
    mem[4006] = 'd188;
    mem[4007] = 'd752;
    mem[4008] = 'd156;
    mem[4009] = 'd736;
    mem[4010] = 'd116;
    mem[4011] = 'd720;
    mem[4012] = 'd92;
    mem[4013] = 'd696;
    mem[4014] = 'd80;
    mem[4015] = 'd668;
    mem[4016] = 'd68;
    mem[4017] = 'd628;
    mem[4018] = 'd44;
    mem[4019] = 'd556;
    mem[4020] = 'd20;
    mem[4021] = 'd464;
    mem[4022] = 'd744;
    mem[4023] = 'd848;
    mem[4024] = 'd1020;
    mem[4025] = 'd1020;
    mem[4026] = 'd1020;
    mem[4027] = 'd1020;
    mem[4028] = 'd1020;
    mem[4029] = 'd1020;
    mem[4030] = 'd1020;
    mem[4031] = 'd1020;
    mem[4032] = 'd876;
    mem[4033] = 'd956;
    mem[4034] = 'd456;
    mem[4035] = 'd836;
    mem[4036] = 'd556;
    mem[4037] = 'd892;
    mem[4038] = 'd624;
    mem[4039] = 'd940;
    mem[4040] = 'd668;
    mem[4041] = 'd980;
    mem[4042] = 'd700;
    mem[4043] = 'd1008;
    mem[4044] = 'd716;
    mem[4045] = 'd1016;
    mem[4046] = 'd736;
    mem[4047] = 'd1020;
    mem[4048] = 'd752;
    mem[4049] = 'd1020;
    mem[4050] = 'd712;
    mem[4051] = 'd912;
    mem[4052] = 'd332;
    mem[4053] = 'd552;
    mem[4054] = 'd252;
    mem[4055] = 'd476;
    mem[4056] = 'd288;
    mem[4057] = 'd520;
    mem[4058] = 'd420;
    mem[4059] = 'd668;
    mem[4060] = 'd548;
    mem[4061] = 'd804;
    mem[4062] = 'd640;
    mem[4063] = 'd892;
    mem[4064] = 'd676;
    mem[4065] = 'd928;
    mem[4066] = 'd672;
    mem[4067] = 'd924;
    mem[4068] = 'd628;
    mem[4069] = 'd880;
    mem[4070] = 'd536;
    mem[4071] = 'd788;
    mem[4072] = 'd404;
    mem[4073] = 'd652;
    mem[4074] = 'd288;
    mem[4075] = 'd516;
    mem[4076] = 'd256;
    mem[4077] = 'd480;
    mem[4078] = 'd372;
    mem[4079] = 'd584;
    mem[4080] = 'd752;
    mem[4081] = 'd956;
    mem[4082] = 'd752;
    mem[4083] = 'd1020;
    mem[4084] = 'd736;
    mem[4085] = 'd1020;
    mem[4086] = 'd720;
    mem[4087] = 'd1016;
    mem[4088] = 'd696;
    mem[4089] = 'd1008;
    mem[4090] = 'd668;
    mem[4091] = 'd980;
    mem[4092] = 'd628;
    mem[4093] = 'd948;
    mem[4094] = 'd556;
    mem[4095] = 'd892;
    mem[4096] = 'd464;
    mem[4097] = 'd836;
    mem[4098] = 'd848;
    mem[4099] = 'd952;
    mem[4100] = 'd1020;
    mem[4101] = 'd1020;
    mem[4102] = 'd1020;
    mem[4103] = 'd1020;
    mem[4104] = 'd1020;
    mem[4105] = 'd1020;
    mem[4106] = 'd1020;
    mem[4107] = 'd1020;
    mem[4108] = 'd1020;
    mem[4109] = 'd1020;
    mem[4110] = 'd280;
    mem[4111] = 'd576;
    mem[4112] = 'd28;
    mem[4113] = 'd504;
    mem[4114] = 'd52;
    mem[4115] = 'd580;
    mem[4116] = 'd72;
    mem[4117] = 'd636;
    mem[4118] = 'd84;
    mem[4119] = 'd672;
    mem[4120] = 'd92;
    mem[4121] = 'd696;
    mem[4122] = 'd108;
    mem[4123] = 'd716;
    mem[4124] = 'd144;
    mem[4125] = 'd732;
    mem[4126] = 'd180;
    mem[4127] = 'd748;
    mem[4128] = 'd224;
    mem[4129] = 'd752;
    mem[4130] = 'd112;
    mem[4131] = 'd480;
    mem[4132] = 'd20;
    mem[4133] = 'd308;
    mem[4134] = 'd20;
    mem[4135] = 'd296;
    mem[4136] = 'd16;
    mem[4137] = 'd264;
    mem[4138] = 'd20;
    mem[4139] = 'd248;
    mem[4140] = 'd20;
    mem[4141] = 'd244;
    mem[4142] = 'd20;
    mem[4143] = 'd248;
    mem[4144] = 'd20;
    mem[4145] = 'd252;
    mem[4146] = 'd16;
    mem[4147] = 'd268;
    mem[4148] = 'd20;
    mem[4149] = 'd300;
    mem[4150] = 'd28;
    mem[4151] = 'd328;
    mem[4152] = 'd136;
    mem[4153] = 'd532;
    mem[4154] = 'd224;
    mem[4155] = 'd768;
    mem[4156] = 'd176;
    mem[4157] = 'd748;
    mem[4158] = 'd144;
    mem[4159] = 'd732;
    mem[4160] = 'd112;
    mem[4161] = 'd716;
    mem[4162] = 'd92;
    mem[4163] = 'd696;
    mem[4164] = 'd84;
    mem[4165] = 'd676;
    mem[4166] = 'd76;
    mem[4167] = 'd640;
    mem[4168] = 'd56;
    mem[4169] = 'd588;
    mem[4170] = 'd32;
    mem[4171] = 'd508;
    mem[4172] = 'd256;
    mem[4173] = 'd564;
    mem[4174] = 'd1008;
    mem[4175] = 'd1012;
    mem[4176] = 'd1020;
    mem[4177] = 'd1020;
    mem[4178] = 'd1020;
    mem[4179] = 'd1020;
    mem[4180] = 'd1020;
    mem[4181] = 'd1020;
    mem[4182] = 'd1020;
    mem[4183] = 'd1020;
    mem[4184] = 'd1020;
    mem[4185] = 'd1020;
    mem[4186] = 'd576;
    mem[4187] = 'd856;
    mem[4188] = 'd504;
    mem[4189] = 'd856;
    mem[4190] = 'd580;
    mem[4191] = 'd904;
    mem[4192] = 'd636;
    mem[4193] = 'd952;
    mem[4194] = 'd672;
    mem[4195] = 'd984;
    mem[4196] = 'd696;
    mem[4197] = 'd1004;
    mem[4198] = 'd716;
    mem[4199] = 'd1020;
    mem[4200] = 'd732;
    mem[4201] = 'd1020;
    mem[4202] = 'd748;
    mem[4203] = 'd1020;
    mem[4204] = 'd752;
    mem[4205] = 'd956;
    mem[4206] = 'd480;
    mem[4207] = 'd680;
    mem[4208] = 'd308;
    mem[4209] = 'd544;
    mem[4210] = 'd296;
    mem[4211] = 'd528;
    mem[4212] = 'd264;
    mem[4213] = 'd488;
    mem[4214] = 'd248;
    mem[4215] = 'd468;
    mem[4216] = 'd244;
    mem[4217] = 'd468;
    mem[4218] = 'd248;
    mem[4219] = 'd468;
    mem[4220] = 'd252;
    mem[4221] = 'd472;
    mem[4222] = 'd268;
    mem[4223] = 'd496;
    mem[4224] = 'd300;
    mem[4225] = 'd528;
    mem[4226] = 'd328;
    mem[4227] = 'd560;
    mem[4228] = 'd532;
    mem[4229] = 'd728;
    mem[4230] = 'd768;
    mem[4231] = 'd976;
    mem[4232] = 'd748;
    mem[4233] = 'd1020;
    mem[4234] = 'd732;
    mem[4235] = 'd1020;
    mem[4236] = 'd716;
    mem[4237] = 'd1020;
    mem[4238] = 'd696;
    mem[4239] = 'd1008;
    mem[4240] = 'd676;
    mem[4241] = 'd984;
    mem[4242] = 'd640;
    mem[4243] = 'd956;
    mem[4244] = 'd588;
    mem[4245] = 'd912;
    mem[4246] = 'd508;
    mem[4247] = 'd860;
    mem[4248] = 'd564;
    mem[4249] = 'd856;
    mem[4250] = 'd1012;
    mem[4251] = 'd1012;
    mem[4252] = 'd1020;
    mem[4253] = 'd1020;
    mem[4254] = 'd1020;
    mem[4255] = 'd1020;
    mem[4256] = 'd1020;
    mem[4257] = 'd1020;
    mem[4258] = 'd1020;
    mem[4259] = 'd1020;
    mem[4260] = 'd1020;
    mem[4261] = 'd1020;
    mem[4262] = 'd848;
    mem[4263] = 'd912;
    mem[4264] = 'd24;
    mem[4265] = 'd456;
    mem[4266] = 'd36;
    mem[4267] = 'd528;
    mem[4268] = 'd60;
    mem[4269] = 'd596;
    mem[4270] = 'd76;
    mem[4271] = 'd640;
    mem[4272] = 'd88;
    mem[4273] = 'd672;
    mem[4274] = 'd92;
    mem[4275] = 'd692;
    mem[4276] = 'd100;
    mem[4277] = 'd708;
    mem[4278] = 'd124;
    mem[4279] = 'd724;
    mem[4280] = 'd152;
    mem[4281] = 'd736;
    mem[4282] = 'd200;
    mem[4283] = 'd768;
    mem[4284] = 'd204;
    mem[4285] = 'd708;
    mem[4286] = 'd132;
    mem[4287] = 'd532;
    mem[4288] = 'd60;
    mem[4289] = 'd400;
    mem[4290] = 'd32;
    mem[4291] = 'd352;
    mem[4292] = 'd24;
    mem[4293] = 'd344;
    mem[4294] = 'd28;
    mem[4295] = 'd344;
    mem[4296] = 'd36;
    mem[4297] = 'd364;
    mem[4298] = 'd72;
    mem[4299] = 'd420;
    mem[4300] = 'd140;
    mem[4301] = 'd556;
    mem[4302] = 'd204;
    mem[4303] = 'd716;
    mem[4304] = 'd192;
    mem[4305] = 'd764;
    mem[4306] = 'd156;
    mem[4307] = 'd736;
    mem[4308] = 'd128;
    mem[4309] = 'd724;
    mem[4310] = 'd100;
    mem[4311] = 'd708;
    mem[4312] = 'd92;
    mem[4313] = 'd692;
    mem[4314] = 'd88;
    mem[4315] = 'd672;
    mem[4316] = 'd80;
    mem[4317] = 'd644;
    mem[4318] = 'd64;
    mem[4319] = 'd600;
    mem[4320] = 'd40;
    mem[4321] = 'd532;
    mem[4322] = 'd52;
    mem[4323] = 'd472;
    mem[4324] = 'd796;
    mem[4325] = 'd880;
    mem[4326] = 'd1020;
    mem[4327] = 'd1020;
    mem[4328] = 'd1020;
    mem[4329] = 'd1020;
    mem[4330] = 'd1020;
    mem[4331] = 'd1020;
    mem[4332] = 'd1020;
    mem[4333] = 'd1020;
    mem[4334] = 'd1020;
    mem[4335] = 'd1020;
    mem[4336] = 'd1020;
    mem[4337] = 'd1020;
    mem[4338] = 'd912;
    mem[4339] = 'd972;
    mem[4340] = 'd456;
    mem[4341] = 'd828;
    mem[4342] = 'd528;
    mem[4343] = 'd868;
    mem[4344] = 'd596;
    mem[4345] = 'd916;
    mem[4346] = 'd640;
    mem[4347] = 'd956;
    mem[4348] = 'd672;
    mem[4349] = 'd984;
    mem[4350] = 'd692;
    mem[4351] = 'd1004;
    mem[4352] = 'd708;
    mem[4353] = 'd1016;
    mem[4354] = 'd724;
    mem[4355] = 'd1020;
    mem[4356] = 'd736;
    mem[4357] = 'd1020;
    mem[4358] = 'd768;
    mem[4359] = 'd1016;
    mem[4360] = 'd708;
    mem[4361] = 'd896;
    mem[4362] = 'd532;
    mem[4363] = 'd728;
    mem[4364] = 'd400;
    mem[4365] = 'd624;
    mem[4366] = 'd352;
    mem[4367] = 'd584;
    mem[4368] = 'd344;
    mem[4369] = 'd576;
    mem[4370] = 'd344;
    mem[4371] = 'd580;
    mem[4372] = 'd364;
    mem[4373] = 'd596;
    mem[4374] = 'd420;
    mem[4375] = 'd640;
    mem[4376] = 'd556;
    mem[4377] = 'd752;
    mem[4378] = 'd716;
    mem[4379] = 'd916;
    mem[4380] = 'd764;
    mem[4381] = 'd1020;
    mem[4382] = 'd736;
    mem[4383] = 'd1020;
    mem[4384] = 'd724;
    mem[4385] = 'd1020;
    mem[4386] = 'd708;
    mem[4387] = 'd1016;
    mem[4388] = 'd692;
    mem[4389] = 'd1008;
    mem[4390] = 'd672;
    mem[4391] = 'd988;
    mem[4392] = 'd644;
    mem[4393] = 'd956;
    mem[4394] = 'd600;
    mem[4395] = 'd920;
    mem[4396] = 'd532;
    mem[4397] = 'd872;
    mem[4398] = 'd472;
    mem[4399] = 'd836;
    mem[4400] = 'd880;
    mem[4401] = 'd964;
    mem[4402] = 'd1020;
    mem[4403] = 'd1020;
    mem[4404] = 'd1020;
    mem[4405] = 'd1020;
    mem[4406] = 'd1020;
    mem[4407] = 'd1020;
    mem[4408] = 'd1020;
    mem[4409] = 'd1020;
    mem[4410] = 'd1020;
    mem[4411] = 'd1020;
    mem[4412] = 'd1020;
    mem[4413] = 'd1020;
    mem[4414] = 'd1016;
    mem[4415] = 'd1020;
    mem[4416] = 'd424;
    mem[4417] = 'd668;
    mem[4418] = 'd20;
    mem[4419] = 'd476;
    mem[4420] = 'd40;
    mem[4421] = 'd540;
    mem[4422] = 'd60;
    mem[4423] = 'd600;
    mem[4424] = 'd80;
    mem[4425] = 'd640;
    mem[4426] = 'd88;
    mem[4427] = 'd664;
    mem[4428] = 'd92;
    mem[4429] = 'd684;
    mem[4430] = 'd96;
    mem[4431] = 'd700;
    mem[4432] = 'd108;
    mem[4433] = 'd712;
    mem[4434] = 'd124;
    mem[4435] = 'd720;
    mem[4436] = 'd144;
    mem[4437] = 'd732;
    mem[4438] = 'd176;
    mem[4439] = 'd752;
    mem[4440] = 'd208;
    mem[4441] = 'd780;
    mem[4442] = 'd216;
    mem[4443] = 'd776;
    mem[4444] = 'd212;
    mem[4445] = 'd756;
    mem[4446] = 'd216;
    mem[4447] = 'd756;
    mem[4448] = 'd212;
    mem[4449] = 'd768;
    mem[4450] = 'd204;
    mem[4451] = 'd776;
    mem[4452] = 'd172;
    mem[4453] = 'd752;
    mem[4454] = 'd144;
    mem[4455] = 'd732;
    mem[4456] = 'd124;
    mem[4457] = 'd720;
    mem[4458] = 'd112;
    mem[4459] = 'd712;
    mem[4460] = 'd100;
    mem[4461] = 'd700;
    mem[4462] = 'd92;
    mem[4463] = 'd684;
    mem[4464] = 'd88;
    mem[4465] = 'd668;
    mem[4466] = 'd80;
    mem[4467] = 'd640;
    mem[4468] = 'd64;
    mem[4469] = 'd604;
    mem[4470] = 'd44;
    mem[4471] = 'd548;
    mem[4472] = 'd20;
    mem[4473] = 'd480;
    mem[4474] = 'd408;
    mem[4475] = 'd660;
    mem[4476] = 'd1016;
    mem[4477] = 'd1020;
    mem[4478] = 'd1020;
    mem[4479] = 'd1020;
    mem[4480] = 'd1020;
    mem[4481] = 'd1020;
    mem[4482] = 'd1020;
    mem[4483] = 'd1020;
    mem[4484] = 'd1020;
    mem[4485] = 'd1020;
    mem[4486] = 'd1020;
    mem[4487] = 'd1020;
    mem[4488] = 'd1020;
    mem[4489] = 'd1020;
    mem[4490] = 'd1020;
    mem[4491] = 'd1020;
    mem[4492] = 'd668;
    mem[4493] = 'd896;
    mem[4494] = 'd476;
    mem[4495] = 'd844;
    mem[4496] = 'd540;
    mem[4497] = 'd876;
    mem[4498] = 'd600;
    mem[4499] = 'd920;
    mem[4500] = 'd640;
    mem[4501] = 'd956;
    mem[4502] = 'd664;
    mem[4503] = 'd980;
    mem[4504] = 'd684;
    mem[4505] = 'd996;
    mem[4506] = 'd700;
    mem[4507] = 'd1012;
    mem[4508] = 'd712;
    mem[4509] = 'd1020;
    mem[4510] = 'd720;
    mem[4511] = 'd1020;
    mem[4512] = 'd732;
    mem[4513] = 'd1020;
    mem[4514] = 'd752;
    mem[4515] = 'd1020;
    mem[4516] = 'd780;
    mem[4517] = 'd1012;
    mem[4518] = 'd776;
    mem[4519] = 'd984;
    mem[4520] = 'd756;
    mem[4521] = 'd960;
    mem[4522] = 'd756;
    mem[4523] = 'd960;
    mem[4524] = 'd768;
    mem[4525] = 'd976;
    mem[4526] = 'd776;
    mem[4527] = 'd1012;
    mem[4528] = 'd752;
    mem[4529] = 'd1020;
    mem[4530] = 'd732;
    mem[4531] = 'd1020;
    mem[4532] = 'd720;
    mem[4533] = 'd1020;
    mem[4534] = 'd712;
    mem[4535] = 'd1020;
    mem[4536] = 'd700;
    mem[4537] = 'd1012;
    mem[4538] = 'd684;
    mem[4539] = 'd1000;
    mem[4540] = 'd668;
    mem[4541] = 'd984;
    mem[4542] = 'd640;
    mem[4543] = 'd956;
    mem[4544] = 'd604;
    mem[4545] = 'd924;
    mem[4546] = 'd548;
    mem[4547] = 'd880;
    mem[4548] = 'd480;
    mem[4549] = 'd844;
    mem[4550] = 'd660;
    mem[4551] = 'd892;
    mem[4552] = 'd1020;
    mem[4553] = 'd1020;
    mem[4554] = 'd1020;
    mem[4555] = 'd1020;
    mem[4556] = 'd1020;
    mem[4557] = 'd1020;
    mem[4558] = 'd1020;
    mem[4559] = 'd1020;
    mem[4560] = 'd1020;
    mem[4561] = 'd1020;
    mem[4562] = 'd1020;
    mem[4563] = 'd1020;
    mem[4564] = 'd1020;
    mem[4565] = 'd1020;
    mem[4566] = 'd1016;
    mem[4567] = 'd1020;
    mem[4568] = 'd948;
    mem[4569] = 'd976;
    mem[4570] = 'd220;
    mem[4571] = 'd540;
    mem[4572] = 'd24;
    mem[4573] = 'd488;
    mem[4574] = 'd44;
    mem[4575] = 'd548;
    mem[4576] = 'd60;
    mem[4577] = 'd596;
    mem[4578] = 'd76;
    mem[4579] = 'd632;
    mem[4580] = 'd84;
    mem[4581] = 'd656;
    mem[4582] = 'd88;
    mem[4583] = 'd672;
    mem[4584] = 'd92;
    mem[4585] = 'd688;
    mem[4586] = 'd96;
    mem[4587] = 'd696;
    mem[4588] = 'd104;
    mem[4589] = 'd704;
    mem[4590] = 'd116;
    mem[4591] = 'd712;
    mem[4592] = 'd128;
    mem[4593] = 'd716;
    mem[4594] = 'd132;
    mem[4595] = 'd716;
    mem[4596] = 'd132;
    mem[4597] = 'd720;
    mem[4598] = 'd132;
    mem[4599] = 'd716;
    mem[4600] = 'd132;
    mem[4601] = 'd716;
    mem[4602] = 'd128;
    mem[4603] = 'd716;
    mem[4604] = 'd120;
    mem[4605] = 'd712;
    mem[4606] = 'd104;
    mem[4607] = 'd704;
    mem[4608] = 'd92;
    mem[4609] = 'd696;
    mem[4610] = 'd92;
    mem[4611] = 'd688;
    mem[4612] = 'd88;
    mem[4613] = 'd676;
    mem[4614] = 'd88;
    mem[4615] = 'd660;
    mem[4616] = 'd80;
    mem[4617] = 'd636;
    mem[4618] = 'd68;
    mem[4619] = 'd600;
    mem[4620] = 'd48;
    mem[4621] = 'd552;
    mem[4622] = 'd24;
    mem[4623] = 'd492;
    mem[4624] = 'd192;
    mem[4625] = 'd520;
    mem[4626] = 'd936;
    mem[4627] = 'd964;
    mem[4628] = 'd1016;
    mem[4629] = 'd1020;
    mem[4630] = 'd1020;
    mem[4631] = 'd1020;
    mem[4632] = 'd1020;
    mem[4633] = 'd1020;
    mem[4634] = 'd1020;
    mem[4635] = 'd1020;
    mem[4636] = 'd1020;
    mem[4637] = 'd1020;
    mem[4638] = 'd1020;
    mem[4639] = 'd1020;
    mem[4640] = 'd1020;
    mem[4641] = 'd1020;
    mem[4642] = 'd1020;
    mem[4643] = 'd1020;
    mem[4644] = 'd976;
    mem[4645] = 'd1000;
    mem[4646] = 'd540;
    mem[4647] = 'd844;
    mem[4648] = 'd488;
    mem[4649] = 'd848;
    mem[4650] = 'd548;
    mem[4651] = 'd880;
    mem[4652] = 'd596;
    mem[4653] = 'd916;
    mem[4654] = 'd632;
    mem[4655] = 'd952;
    mem[4656] = 'd656;
    mem[4657] = 'd972;
    mem[4658] = 'd672;
    mem[4659] = 'd992;
    mem[4660] = 'd688;
    mem[4661] = 'd1004;
    mem[4662] = 'd696;
    mem[4663] = 'd1016;
    mem[4664] = 'd704;
    mem[4665] = 'd1020;
    mem[4666] = 'd712;
    mem[4667] = 'd1020;
    mem[4668] = 'd716;
    mem[4669] = 'd1020;
    mem[4670] = 'd716;
    mem[4671] = 'd1020;
    mem[4672] = 'd720;
    mem[4673] = 'd1020;
    mem[4674] = 'd716;
    mem[4675] = 'd1020;
    mem[4676] = 'd716;
    mem[4677] = 'd1020;
    mem[4678] = 'd716;
    mem[4679] = 'd1020;
    mem[4680] = 'd712;
    mem[4681] = 'd1020;
    mem[4682] = 'd704;
    mem[4683] = 'd1020;
    mem[4684] = 'd696;
    mem[4685] = 'd1016;
    mem[4686] = 'd688;
    mem[4687] = 'd1008;
    mem[4688] = 'd676;
    mem[4689] = 'd992;
    mem[4690] = 'd660;
    mem[4691] = 'd976;
    mem[4692] = 'd636;
    mem[4693] = 'd952;
    mem[4694] = 'd600;
    mem[4695] = 'd920;
    mem[4696] = 'd552;
    mem[4697] = 'd884;
    mem[4698] = 'd492;
    mem[4699] = 'd852;
    mem[4700] = 'd520;
    mem[4701] = 'd836;
    mem[4702] = 'd964;
    mem[4703] = 'd996;
    mem[4704] = 'd1020;
    mem[4705] = 'd1020;
    mem[4706] = 'd1020;
    mem[4707] = 'd1020;
    mem[4708] = 'd1020;
    mem[4709] = 'd1020;
    mem[4710] = 'd1020;
    mem[4711] = 'd1020;
    mem[4712] = 'd1020;
    mem[4713] = 'd1020;
    mem[4714] = 'd1020;
    mem[4715] = 'd1020;
    mem[4716] = 'd1020;
    mem[4717] = 'd1020;
    mem[4718] = 'd1020;
    mem[4719] = 'd1020;
    mem[4720] = 'd1016;
    mem[4721] = 'd1020;
    mem[4722] = 'd900;
    mem[4723] = 'd944;
    mem[4724] = 'd168;
    mem[4725] = 'd504;
    mem[4726] = 'd24;
    mem[4727] = 'd488;
    mem[4728] = 'd40;
    mem[4729] = 'd540;
    mem[4730] = 'd56;
    mem[4731] = 'd584;
    mem[4732] = 'd72;
    mem[4733] = 'd620;
    mem[4734] = 'd80;
    mem[4735] = 'd644;
    mem[4736] = 'd88;
    mem[4737] = 'd660;
    mem[4738] = 'd88;
    mem[4739] = 'd672;
    mem[4740] = 'd92;
    mem[4741] = 'd680;
    mem[4742] = 'd92;
    mem[4743] = 'd688;
    mem[4744] = 'd92;
    mem[4745] = 'd692;
    mem[4746] = 'd96;
    mem[4747] = 'd692;
    mem[4748] = 'd96;
    mem[4749] = 'd692;
    mem[4750] = 'd100;
    mem[4751] = 'd696;
    mem[4752] = 'd96;
    mem[4753] = 'd692;
    mem[4754] = 'd92;
    mem[4755] = 'd692;
    mem[4756] = 'd92;
    mem[4757] = 'd684;
    mem[4758] = 'd92;
    mem[4759] = 'd680;
    mem[4760] = 'd88;
    mem[4761] = 'd676;
    mem[4762] = 'd88;
    mem[4763] = 'd664;
    mem[4764] = 'd84;
    mem[4765] = 'd648;
    mem[4766] = 'd76;
    mem[4767] = 'd624;
    mem[4768] = 'd60;
    mem[4769] = 'd588;
    mem[4770] = 'd44;
    mem[4771] = 'd548;
    mem[4772] = 'd24;
    mem[4773] = 'd492;
    mem[4774] = 'd144;
    mem[4775] = 'd496;
    mem[4776] = 'd892;
    mem[4777] = 'd940;
    mem[4778] = 'd1016;
    mem[4779] = 'd1020;
    mem[4780] = 'd1020;
    mem[4781] = 'd1020;
    mem[4782] = 'd1020;
    mem[4783] = 'd1020;
    mem[4784] = 'd1020;
    mem[4785] = 'd1020;
    mem[4786] = 'd1020;
    mem[4787] = 'd1020;
    mem[4788] = 'd1020;
    mem[4789] = 'd1020;
    mem[4790] = 'd1020;
    mem[4791] = 'd1020;
    mem[4792] = 'd1020;
    mem[4793] = 'd1020;
    mem[4794] = 'd1020;
    mem[4795] = 'd1020;
    mem[4796] = 'd1020;
    mem[4797] = 'd1020;
    mem[4798] = 'd944;
    mem[4799] = 'd988;
    mem[4800] = 'd504;
    mem[4801] = 'd824;
    mem[4802] = 'd488;
    mem[4803] = 'd852;
    mem[4804] = 'd540;
    mem[4805] = 'd880;
    mem[4806] = 'd584;
    mem[4807] = 'd908;
    mem[4808] = 'd620;
    mem[4809] = 'd940;
    mem[4810] = 'd644;
    mem[4811] = 'd960;
    mem[4812] = 'd660;
    mem[4813] = 'd980;
    mem[4814] = 'd672;
    mem[4815] = 'd996;
    mem[4816] = 'd680;
    mem[4817] = 'd1004;
    mem[4818] = 'd688;
    mem[4819] = 'd1012;
    mem[4820] = 'd692;
    mem[4821] = 'd1016;
    mem[4822] = 'd692;
    mem[4823] = 'd1016;
    mem[4824] = 'd692;
    mem[4825] = 'd1016;
    mem[4826] = 'd696;
    mem[4827] = 'd1016;
    mem[4828] = 'd692;
    mem[4829] = 'd1016;
    mem[4830] = 'd692;
    mem[4831] = 'd1016;
    mem[4832] = 'd684;
    mem[4833] = 'd1012;
    mem[4834] = 'd680;
    mem[4835] = 'd1004;
    mem[4836] = 'd676;
    mem[4837] = 'd996;
    mem[4838] = 'd664;
    mem[4839] = 'd984;
    mem[4840] = 'd648;
    mem[4841] = 'd968;
    mem[4842] = 'd624;
    mem[4843] = 'd940;
    mem[4844] = 'd588;
    mem[4845] = 'd912;
    mem[4846] = 'd548;
    mem[4847] = 'd884;
    mem[4848] = 'd492;
    mem[4849] = 'd852;
    mem[4850] = 'd496;
    mem[4851] = 'd828;
    mem[4852] = 'd940;
    mem[4853] = 'd988;
    mem[4854] = 'd1020;
    mem[4855] = 'd1020;
    mem[4856] = 'd1020;
    mem[4857] = 'd1020;
    mem[4858] = 'd1020;
    mem[4859] = 'd1020;
    mem[4860] = 'd1020;
    mem[4861] = 'd1020;
    mem[4862] = 'd1020;
    mem[4863] = 'd1020;
    mem[4864] = 'd1020;
    mem[4865] = 'd1020;
    mem[4866] = 'd1020;
    mem[4867] = 'd1020;
    mem[4868] = 'd1020;
    mem[4869] = 'd1020;
    mem[4870] = 'd1020;
    mem[4871] = 'd1020;
    mem[4872] = 'd1016;
    mem[4873] = 'd1020;
    mem[4874] = 'd1012;
    mem[4875] = 'd1020;
    mem[4876] = 'd896;
    mem[4877] = 'd940;
    mem[4878] = 'd220;
    mem[4879] = 'd540;
    mem[4880] = 'd20;
    mem[4881] = 'd476;
    mem[4882] = 'd36;
    mem[4883] = 'd528;
    mem[4884] = 'd52;
    mem[4885] = 'd572;
    mem[4886] = 'd64;
    mem[4887] = 'd600;
    mem[4888] = 'd72;
    mem[4889] = 'd624;
    mem[4890] = 'd80;
    mem[4891] = 'd640;
    mem[4892] = 'd84;
    mem[4893] = 'd656;
    mem[4894] = 'd88;
    mem[4895] = 'd664;
    mem[4896] = 'd88;
    mem[4897] = 'd668;
    mem[4898] = 'd92;
    mem[4899] = 'd672;
    mem[4900] = 'd88;
    mem[4901] = 'd672;
    mem[4902] = 'd88;
    mem[4903] = 'd672;
    mem[4904] = 'd88;
    mem[4905] = 'd672;
    mem[4906] = 'd88;
    mem[4907] = 'd668;
    mem[4908] = 'd88;
    mem[4909] = 'd664;
    mem[4910] = 'd84;
    mem[4911] = 'd656;
    mem[4912] = 'd80;
    mem[4913] = 'd644;
    mem[4914] = 'd72;
    mem[4915] = 'd628;
    mem[4916] = 'd64;
    mem[4917] = 'd604;
    mem[4918] = 'd56;
    mem[4919] = 'd572;
    mem[4920] = 'd36;
    mem[4921] = 'd532;
    mem[4922] = 'd24;
    mem[4923] = 'd480;
    mem[4924] = 'd196;
    mem[4925] = 'd520;
    mem[4926] = 'd892;
    mem[4927] = 'd940;
    mem[4928] = 'd1012;
    mem[4929] = 'd1016;
    mem[4930] = 'd1016;
    mem[4931] = 'd1020;
    mem[4932] = 'd1020;
    mem[4933] = 'd1020;
    mem[4934] = 'd1020;
    mem[4935] = 'd1020;
    mem[4936] = 'd1020;
    mem[4937] = 'd1020;
    mem[4938] = 'd1020;
    mem[4939] = 'd1020;
    mem[4940] = 'd1020;
    mem[4941] = 'd1020;
    mem[4942] = 'd1020;
    mem[4943] = 'd1020;
    mem[4944] = 'd1020;
    mem[4945] = 'd1020;
    mem[4946] = 'd1020;
    mem[4947] = 'd1020;
    mem[4948] = 'd1020;
    mem[4949] = 'd1020;
    mem[4950] = 'd1020;
    mem[4951] = 'd1020;
    mem[4952] = 'd940;
    mem[4953] = 'd988;
    mem[4954] = 'd540;
    mem[4955] = 'd840;
    mem[4956] = 'd476;
    mem[4957] = 'd844;
    mem[4958] = 'd528;
    mem[4959] = 'd876;
    mem[4960] = 'd572;
    mem[4961] = 'd900;
    mem[4962] = 'd600;
    mem[4963] = 'd924;
    mem[4964] = 'd624;
    mem[4965] = 'd948;
    mem[4966] = 'd640;
    mem[4967] = 'd964;
    mem[4968] = 'd656;
    mem[4969] = 'd980;
    mem[4970] = 'd664;
    mem[4971] = 'd988;
    mem[4972] = 'd668;
    mem[4973] = 'd996;
    mem[4974] = 'd672;
    mem[4975] = 'd996;
    mem[4976] = 'd672;
    mem[4977] = 'd1000;
    mem[4978] = 'd672;
    mem[4979] = 'd1000;
    mem[4980] = 'd672;
    mem[4981] = 'd996;
    mem[4982] = 'd668;
    mem[4983] = 'd996;
    mem[4984] = 'd664;
    mem[4985] = 'd988;
    mem[4986] = 'd656;
    mem[4987] = 'd980;
    mem[4988] = 'd644;
    mem[4989] = 'd964;
    mem[4990] = 'd628;
    mem[4991] = 'd948;
    mem[4992] = 'd604;
    mem[4993] = 'd928;
    mem[4994] = 'd572;
    mem[4995] = 'd904;
    mem[4996] = 'd532;
    mem[4997] = 'd880;
    mem[4998] = 'd480;
    mem[4999] = 'd848;
    mem[5000] = 'd520;
    mem[5001] = 'd832;
    mem[5002] = 'd940;
    mem[5003] = 'd988;
    mem[5004] = 'd1016;
    mem[5005] = 'd1020;
    mem[5006] = 'd1020;
    mem[5007] = 'd1020;
    mem[5008] = 'd1020;
    mem[5009] = 'd1020;
    mem[5010] = 'd1020;
    mem[5011] = 'd1020;
    mem[5012] = 'd1020;
    mem[5013] = 'd1020;
    mem[5014] = 'd1020;
    mem[5015] = 'd1020;
    mem[5016] = 'd1020;
    mem[5017] = 'd1020;
    mem[5018] = 'd1020;
    mem[5019] = 'd1020;
    mem[5020] = 'd1020;
    mem[5021] = 'd1020;
    mem[5022] = 'd1020;
    mem[5023] = 'd1020;
    mem[5024] = 'd1020;
    mem[5025] = 'd1020;
    mem[5026] = 'd1016;
    mem[5027] = 'd1020;
    mem[5028] = 'd1012;
    mem[5029] = 'd1020;
    mem[5030] = 'd944;
    mem[5031] = 'd976;
    mem[5032] = 'd416;
    mem[5033] = 'd664;
    mem[5034] = 'd24;
    mem[5035] = 'd456;
    mem[5036] = 'd28;
    mem[5037] = 'd504;
    mem[5038] = 'd40;
    mem[5039] = 'd544;
    mem[5040] = 'd52;
    mem[5041] = 'd576;
    mem[5042] = 'd60;
    mem[5043] = 'd596;
    mem[5044] = 'd68;
    mem[5045] = 'd616;
    mem[5046] = 'd72;
    mem[5047] = 'd628;
    mem[5048] = 'd76;
    mem[5049] = 'd636;
    mem[5050] = 'd80;
    mem[5051] = 'd644;
    mem[5052] = 'd80;
    mem[5053] = 'd644;
    mem[5054] = 'd80;
    mem[5055] = 'd644;
    mem[5056] = 'd80;
    mem[5057] = 'd640;
    mem[5058] = 'd76;
    mem[5059] = 'd636;
    mem[5060] = 'd72;
    mem[5061] = 'd628;
    mem[5062] = 'd68;
    mem[5063] = 'd620;
    mem[5064] = 'd60;
    mem[5065] = 'd600;
    mem[5066] = 'd52;
    mem[5067] = 'd580;
    mem[5068] = 'd44;
    mem[5069] = 'd548;
    mem[5070] = 'd32;
    mem[5071] = 'd508;
    mem[5072] = 'd24;
    mem[5073] = 'd456;
    mem[5074] = 'd388;
    mem[5075] = 'd648;
    mem[5076] = 'd932;
    mem[5077] = 'd968;
    mem[5078] = 'd1012;
    mem[5079] = 'd1016;
    mem[5080] = 'd1016;
    mem[5081] = 'd1020;
    mem[5082] = 'd1020;
    mem[5083] = 'd1020;
    mem[5084] = 'd1020;
    mem[5085] = 'd1020;
    mem[5086] = 'd1020;
    mem[5087] = 'd1020;
    mem[5088] = 'd1020;
    mem[5089] = 'd1020;
    mem[5090] = 'd1020;
    mem[5091] = 'd1020;
    mem[5092] = 'd1020;
    mem[5093] = 'd1020;
    mem[5094] = 'd1020;
    mem[5095] = 'd1020;
    mem[5096] = 'd1020;
    mem[5097] = 'd1020;
    mem[5098] = 'd1020;
    mem[5099] = 'd1020;
    mem[5100] = 'd1020;
    mem[5101] = 'd1020;
    mem[5102] = 'd1020;
    mem[5103] = 'd1020;
    mem[5104] = 'd1020;
    mem[5105] = 'd1020;
    mem[5106] = 'd976;
    mem[5107] = 'd1000;
    mem[5108] = 'd664;
    mem[5109] = 'd888;
    mem[5110] = 'd456;
    mem[5111] = 'd824;
    mem[5112] = 'd504;
    mem[5113] = 'd864;
    mem[5114] = 'd544;
    mem[5115] = 'd888;
    mem[5116] = 'd576;
    mem[5117] = 'd908;
    mem[5118] = 'd596;
    mem[5119] = 'd924;
    mem[5120] = 'd616;
    mem[5121] = 'd944;
    mem[5122] = 'd628;
    mem[5123] = 'd952;
    mem[5124] = 'd636;
    mem[5125] = 'd964;
    mem[5126] = 'd644;
    mem[5127] = 'd964;
    mem[5128] = 'd644;
    mem[5129] = 'd968;
    mem[5130] = 'd644;
    mem[5131] = 'd968;
    mem[5132] = 'd640;
    mem[5133] = 'd968;
    mem[5134] = 'd636;
    mem[5135] = 'd964;
    mem[5136] = 'd628;
    mem[5137] = 'd956;
    mem[5138] = 'd620;
    mem[5139] = 'd944;
    mem[5140] = 'd600;
    mem[5141] = 'd928;
    mem[5142] = 'd580;
    mem[5143] = 'd912;
    mem[5144] = 'd548;
    mem[5145] = 'd892;
    mem[5146] = 'd508;
    mem[5147] = 'd868;
    mem[5148] = 'd456;
    mem[5149] = 'd828;
    mem[5150] = 'd648;
    mem[5151] = 'd884;
    mem[5152] = 'd968;
    mem[5153] = 'd1000;
    mem[5154] = 'd1016;
    mem[5155] = 'd1020;
    mem[5156] = 'd1020;
    mem[5157] = 'd1020;
    mem[5158] = 'd1020;
    mem[5159] = 'd1020;
    mem[5160] = 'd1020;
    mem[5161] = 'd1020;
    mem[5162] = 'd1020;
    mem[5163] = 'd1020;
    mem[5164] = 'd1020;
    mem[5165] = 'd1020;
    mem[5166] = 'd1020;
    mem[5167] = 'd1020;
    mem[5168] = 'd1020;
    mem[5169] = 'd1020;
    mem[5170] = 'd1020;
    mem[5171] = 'd1020;
    mem[5172] = 'd1020;
    mem[5173] = 'd1020;
    mem[5174] = 'd1020;
    mem[5175] = 'd1020;
    mem[5176] = 'd1020;
    mem[5177] = 'd1020;
    mem[5178] = 'd1020;
    mem[5179] = 'd1020;
    mem[5180] = 'd1016;
    mem[5181] = 'd1020;
    mem[5182] = 'd1012;
    mem[5183] = 'd1020;
    mem[5184] = 'd1004;
    mem[5185] = 'd1012;
    mem[5186] = 'd708;
    mem[5187] = 'd832;
    mem[5188] = 'd180;
    mem[5189] = 'd520;
    mem[5190] = 'd16;
    mem[5191] = 'd460;
    mem[5192] = 'd28;
    mem[5193] = 'd508;
    mem[5194] = 'd40;
    mem[5195] = 'd536;
    mem[5196] = 'd48;
    mem[5197] = 'd560;
    mem[5198] = 'd52;
    mem[5199] = 'd580;
    mem[5200] = 'd56;
    mem[5201] = 'd588;
    mem[5202] = 'd60;
    mem[5203] = 'd596;
    mem[5204] = 'd60;
    mem[5205] = 'd600;
    mem[5206] = 'd60;
    mem[5207] = 'd600;
    mem[5208] = 'd60;
    mem[5209] = 'd600;
    mem[5210] = 'd56;
    mem[5211] = 'd592;
    mem[5212] = 'd52;
    mem[5213] = 'd580;
    mem[5214] = 'd48;
    mem[5215] = 'd564;
    mem[5216] = 'd40;
    mem[5217] = 'd540;
    mem[5218] = 'd28;
    mem[5219] = 'd508;
    mem[5220] = 'd20;
    mem[5221] = 'd464;
    mem[5222] = 'd168;
    mem[5223] = 'd512;
    mem[5224] = 'd680;
    mem[5225] = 'd820;
    mem[5226] = 'd1000;
    mem[5227] = 'd1012;
    mem[5228] = 'd1012;
    mem[5229] = 'd1016;
    mem[5230] = 'd1016;
    mem[5231] = 'd1020;
    mem[5232] = 'd1020;
    mem[5233] = 'd1020;
    mem[5234] = 'd1020;
    mem[5235] = 'd1020;
    mem[5236] = 'd1020;
    mem[5237] = 'd1020;
    mem[5238] = 'd1020;
    mem[5239] = 'd1020;
    mem[5240] = 'd1020;
    mem[5241] = 'd1020;
    mem[5242] = 'd1020;
    mem[5243] = 'd1020;
    mem[5244] = 'd1020;
    mem[5245] = 'd1020;
    mem[5246] = 'd1020;
    mem[5247] = 'd1020;
    mem[5248] = 'd1020;
    mem[5249] = 'd1020;
    mem[5250] = 'd1020;
    mem[5251] = 'd1020;
    mem[5252] = 'd1020;
    mem[5253] = 'd1020;
    mem[5254] = 'd1020;
    mem[5255] = 'd1020;
    mem[5256] = 'd1020;
    mem[5257] = 'd1020;
    mem[5258] = 'd1020;
    mem[5259] = 'd1020;
    mem[5260] = 'd1012;
    mem[5261] = 'd1020;
    mem[5262] = 'd832;
    mem[5263] = 'd944;
    mem[5264] = 'd520;
    mem[5265] = 'd832;
    mem[5266] = 'd460;
    mem[5267] = 'd836;
    mem[5268] = 'd508;
    mem[5269] = 'd868;
    mem[5270] = 'd536;
    mem[5271] = 'd888;
    mem[5272] = 'd560;
    mem[5273] = 'd904;
    mem[5274] = 'd580;
    mem[5275] = 'd912;
    mem[5276] = 'd588;
    mem[5277] = 'd924;
    mem[5278] = 'd596;
    mem[5279] = 'd928;
    mem[5280] = 'd600;
    mem[5281] = 'd932;
    mem[5282] = 'd600;
    mem[5283] = 'd932;
    mem[5284] = 'd600;
    mem[5285] = 'd932;
    mem[5286] = 'd592;
    mem[5287] = 'd924;
    mem[5288] = 'd580;
    mem[5289] = 'd916;
    mem[5290] = 'd564;
    mem[5291] = 'd904;
    mem[5292] = 'd540;
    mem[5293] = 'd888;
    mem[5294] = 'd508;
    mem[5295] = 'd868;
    mem[5296] = 'd464;
    mem[5297] = 'd840;
    mem[5298] = 'd512;
    mem[5299] = 'd832;
    mem[5300] = 'd820;
    mem[5301] = 'd940;
    mem[5302] = 'd1012;
    mem[5303] = 'd1020;
    mem[5304] = 'd1016;
    mem[5305] = 'd1020;
    mem[5306] = 'd1020;
    mem[5307] = 'd1020;
    mem[5308] = 'd1020;
    mem[5309] = 'd1020;
    mem[5310] = 'd1020;
    mem[5311] = 'd1020;
    mem[5312] = 'd1020;
    mem[5313] = 'd1020;
    mem[5314] = 'd1020;
    mem[5315] = 'd1020;
    mem[5316] = 'd1020;
    mem[5317] = 'd1020;
    mem[5318] = 'd1020;
    mem[5319] = 'd1020;
    mem[5320] = 'd1020;
    mem[5321] = 'd1020;
    mem[5322] = 'd1020;
    mem[5323] = 'd1020;
    mem[5324] = 'd1020;
    mem[5325] = 'd1020;
    mem[5326] = 'd1020;
    mem[5327] = 'd1020;
    mem[5328] = 'd1020;
    mem[5329] = 'd1020;
    mem[5330] = 'd1020;
    mem[5331] = 'd1020;
    mem[5332] = 'd1020;
    mem[5333] = 'd1020;
    mem[5334] = 'd1020;
    mem[5335] = 'd1020;
    mem[5336] = 'd1016;
    mem[5337] = 'd1020;
    mem[5338] = 'd1008;
    mem[5339] = 'd1016;
    mem[5340] = 'd968;
    mem[5341] = 'd992;
    mem[5342] = 'd724;
    mem[5343] = 'd840;
    mem[5344] = 'd336;
    mem[5345] = 'd604;
    mem[5346] = 'd68;
    mem[5347] = 'd464;
    mem[5348] = 'd16;
    mem[5349] = 'd468;
    mem[5350] = 'd24;
    mem[5351] = 'd496;
    mem[5352] = 'd28;
    mem[5353] = 'd512;
    mem[5354] = 'd32;
    mem[5355] = 'd524;
    mem[5356] = 'd32;
    mem[5357] = 'd528;
    mem[5358] = 'd32;
    mem[5359] = 'd528;
    mem[5360] = 'd32;
    mem[5361] = 'd524;
    mem[5362] = 'd32;
    mem[5363] = 'd512;
    mem[5364] = 'd24;
    mem[5365] = 'd496;
    mem[5366] = 'd20;
    mem[5367] = 'd472;
    mem[5368] = 'd32;
    mem[5369] = 'd436;
    mem[5370] = 'd328;
    mem[5371] = 'd608;
    mem[5372] = 'd720;
    mem[5373] = 'd836;
    mem[5374] = 'd972;
    mem[5375] = 'd996;
    mem[5376] = 'd1008;
    mem[5377] = 'd1016;
    mem[5378] = 'd1012;
    mem[5379] = 'd1020;
    mem[5380] = 'd1016;
    mem[5381] = 'd1020;
    mem[5382] = 'd1020;
    mem[5383] = 'd1020;
    mem[5384] = 'd1020;
    mem[5385] = 'd1020;
    mem[5386] = 'd1020;
    mem[5387] = 'd1020;
    mem[5388] = 'd1020;
    mem[5389] = 'd1020;
    mem[5390] = 'd1020;
    mem[5391] = 'd1020;
    mem[5392] = 'd1020;
    mem[5393] = 'd1020;
    mem[5394] = 'd1020;
    mem[5395] = 'd1020;
    mem[5396] = 'd1020;
    mem[5397] = 'd1020;
    mem[5398] = 'd1020;
    mem[5399] = 'd1020;
    mem[5400] = 'd1020;
    mem[5401] = 'd1020;
    mem[5402] = 'd1020;
    mem[5403] = 'd1020;
    mem[5404] = 'd1020;
    mem[5405] = 'd1020;
    mem[5406] = 'd1020;
    mem[5407] = 'd1020;
    mem[5408] = 'd1020;
    mem[5409] = 'd1020;
    mem[5410] = 'd1020;
    mem[5411] = 'd1020;
    mem[5412] = 'd1020;
    mem[5413] = 'd1020;
    mem[5414] = 'd1016;
    mem[5415] = 'd1020;
    mem[5416] = 'd992;
    mem[5417] = 'd1008;
    mem[5418] = 'd840;
    mem[5419] = 'd952;
    mem[5420] = 'd604;
    mem[5421] = 'd856;
    mem[5422] = 'd464;
    mem[5423] = 'd816;
    mem[5424] = 'd468;
    mem[5425] = 'd840;
    mem[5426] = 'd496;
    mem[5427] = 'd860;
    mem[5428] = 'd512;
    mem[5429] = 'd872;
    mem[5430] = 'd524;
    mem[5431] = 'd876;
    mem[5432] = 'd528;
    mem[5433] = 'd880;
    mem[5434] = 'd528;
    mem[5435] = 'd880;
    mem[5436] = 'd524;
    mem[5437] = 'd876;
    mem[5438] = 'd512;
    mem[5439] = 'd872;
    mem[5440] = 'd496;
    mem[5441] = 'd860;
    mem[5442] = 'd472;
    mem[5443] = 'd840;
    mem[5444] = 'd436;
    mem[5445] = 'd804;
    mem[5446] = 'd608;
    mem[5447] = 'd860;
    mem[5448] = 'd836;
    mem[5449] = 'd948;
    mem[5450] = 'd996;
    mem[5451] = 'd1012;
    mem[5452] = 'd1016;
    mem[5453] = 'd1020;
    mem[5454] = 'd1020;
    mem[5455] = 'd1020;
    mem[5456] = 'd1020;
    mem[5457] = 'd1020;
    mem[5458] = 'd1020;
    mem[5459] = 'd1020;
    mem[5460] = 'd1020;
    mem[5461] = 'd1020;
    mem[5462] = 'd1020;
    mem[5463] = 'd1020;
    mem[5464] = 'd1020;
    mem[5465] = 'd1020;
    mem[5466] = 'd1020;
    mem[5467] = 'd1020;
    mem[5468] = 'd1020;
    mem[5469] = 'd1020;
    mem[5470] = 'd1020;
    mem[5471] = 'd1020;
    mem[5472] = 'd1020;
    mem[5473] = 'd1020;
    mem[5474] = 'd1020;
    mem[5475] = 'd1020;
    mem[5476] = 'd1020;
    mem[5477] = 'd1020;
    mem[5478] = 'd1020;
    mem[5479] = 'd1020;
    mem[5480] = 'd1020;
    mem[5481] = 'd1020;
    mem[5482] = 'd1020;
    mem[5483] = 'd1020;
    mem[5484] = 'd1020;
    mem[5485] = 'd1020;
    mem[5486] = 'd1020;
    mem[5487] = 'd1020;
    mem[5488] = 'd1020;
    mem[5489] = 'd1020;
    mem[5490] = 'd1016;
    mem[5491] = 'd1020;
    mem[5492] = 'd1012;
    mem[5493] = 'd1016;
    mem[5494] = 'd1012;
    mem[5495] = 'd1016;
    mem[5496] = 'd1008;
    mem[5497] = 'd1016;
    mem[5498] = 'd916;
    mem[5499] = 'd964;
    mem[5500] = 'd652;
    mem[5501] = 'd788;
    mem[5502] = 'd424;
    mem[5503] = 'd652;
    mem[5504] = 'd252;
    mem[5505] = 'd556;
    mem[5506] = 'd148;
    mem[5507] = 'd496;
    mem[5508] = 'd100;
    mem[5509] = 'd472;
    mem[5510] = 'd100;
    mem[5511] = 'd472;
    mem[5512] = 'd144;
    mem[5513] = 'd496;
    mem[5514] = 'd248;
    mem[5515] = 'd552;
    mem[5516] = 'd416;
    mem[5517] = 'd648;
    mem[5518] = 'd652;
    mem[5519] = 'd792;
    mem[5520] = 'd952;
    mem[5521] = 'd984;
    mem[5522] = 'd1004;
    mem[5523] = 'd1016;
    mem[5524] = 'd1012;
    mem[5525] = 'd1016;
    mem[5526] = 'd1016;
    mem[5527] = 'd1020;
    mem[5528] = 'd1016;
    mem[5529] = 'd1020;
    mem[5530] = 'd1020;
    mem[5531] = 'd1020;
    mem[5532] = 'd1020;
    mem[5533] = 'd1020;
    mem[5534] = 'd1020;
    mem[5535] = 'd1020;
    mem[5536] = 'd1020;
    mem[5537] = 'd1020;
    mem[5538] = 'd1020;
    mem[5539] = 'd1020;
    mem[5540] = 'd1020;
    mem[5541] = 'd1020;
    mem[5542] = 'd1020;
    mem[5543] = 'd1020;
    mem[5544] = 'd1020;
    mem[5545] = 'd1020;
    mem[5546] = 'd1020;
    mem[5547] = 'd1020;
    mem[5548] = 'd1020;
    mem[5549] = 'd1020;
    mem[5550] = 'd1020;
    mem[5551] = 'd1020;
    mem[5552] = 'd1020;
    mem[5553] = 'd1020;
    mem[5554] = 'd1020;
    mem[5555] = 'd1020;
    mem[5556] = 'd1020;
    mem[5557] = 'd1020;
    mem[5558] = 'd1020;
    mem[5559] = 'd1020;
    mem[5560] = 'd1020;
    mem[5561] = 'd1020;
    mem[5562] = 'd1020;
    mem[5563] = 'd1020;
    mem[5564] = 'd1020;
    mem[5565] = 'd1020;
    mem[5566] = 'd1020;
    mem[5567] = 'd1020;
    mem[5568] = 'd1016;
    mem[5569] = 'd1020;
    mem[5570] = 'd1016;
    mem[5571] = 'd1020;
    mem[5572] = 'd1016;
    mem[5573] = 'd1020;
    mem[5574] = 'd964;
    mem[5575] = 'd996;
    mem[5576] = 'd788;
    mem[5577] = 'd924;
    mem[5578] = 'd652;
    mem[5579] = 'd868;
    mem[5580] = 'd556;
    mem[5581] = 'd836;
    mem[5582] = 'd496;
    mem[5583] = 'd816;
    mem[5584] = 'd472;
    mem[5585] = 'd808;
    mem[5586] = 'd472;
    mem[5587] = 'd808;
    mem[5588] = 'd496;
    mem[5589] = 'd816;
    mem[5590] = 'd552;
    mem[5591] = 'd836;
    mem[5592] = 'd648;
    mem[5593] = 'd868;
    mem[5594] = 'd792;
    mem[5595] = 'd920;
    mem[5596] = 'd984;
    mem[5597] = 'd1008;
    mem[5598] = 'd1016;
    mem[5599] = 'd1020;
    mem[5600] = 'd1016;
    mem[5601] = 'd1020;
    mem[5602] = 'd1020;
    mem[5603] = 'd1020;
    mem[5604] = 'd1020;
    mem[5605] = 'd1020;
    mem[5606] = 'd1020;
    mem[5607] = 'd1020;
    mem[5608] = 'd1020;
    mem[5609] = 'd1020;
    mem[5610] = 'd1020;
    mem[5611] = 'd1020;
    mem[5612] = 'd1020;
    mem[5613] = 'd1020;
    mem[5614] = 'd1020;
    mem[5615] = 'd1020;
    mem[5616] = 'd1020;
    mem[5617] = 'd1020;
    mem[5618] = 'd1020;
    mem[5619] = 'd1020;
    mem[5620] = 'd1020;
    mem[5621] = 'd1020;
    mem[5622] = 'd1020;
    mem[5623] = 'd1020;
    mem[5624] = 'd1020;
    mem[5625] = 'd1020;
    mem[5626] = 'd1020;
    mem[5627] = 'd1020;
    mem[5628] = 'd1020;
    mem[5629] = 'd1020;
    mem[5630] = 'd1020;
    mem[5631] = 'd1020;
    mem[5632] = 'd1020;
    mem[5633] = 'd1020;
    mem[5634] = 'd1020;
    mem[5635] = 'd1020;
    mem[5636] = 'd1020;
    mem[5637] = 'd1020;
    mem[5638] = 'd1020;
    mem[5639] = 'd1020;
    mem[5640] = 'd1020;
    mem[5641] = 'd1020;
    mem[5642] = 'd1020;
    mem[5643] = 'd1020;
    mem[5644] = 'd1020;
    mem[5645] = 'd1020;
    mem[5646] = 'd1016;
    mem[5647] = 'd1020;
    mem[5648] = 'd1016;
    mem[5649] = 'd1020;
    mem[5650] = 'd1012;
    mem[5651] = 'd1016;
    mem[5652] = 'd1012;
    mem[5653] = 'd1016;
    mem[5654] = 'd1008;
    mem[5655] = 'd1016;
    mem[5656] = 'd1008;
    mem[5657] = 'd1016;
    mem[5658] = 'd1008;
    mem[5659] = 'd1016;
    mem[5660] = 'd1004;
    mem[5661] = 'd1012;
    mem[5662] = 'd1000;
    mem[5663] = 'd1012;
    mem[5664] = 'd1008;
    mem[5665] = 'd1016;
    mem[5666] = 'd1008;
    mem[5667] = 'd1016;
    mem[5668] = 'd1008;
    mem[5669] = 'd1016;
    mem[5670] = 'd1008;
    mem[5671] = 'd1016;
    mem[5672] = 'd1012;
    mem[5673] = 'd1016;
    mem[5674] = 'd1016;
    mem[5675] = 'd1020;
    mem[5676] = 'd1016;
    mem[5677] = 'd1020;
    mem[5678] = 'd1020;
    mem[5679] = 'd1020;
    mem[5680] = 'd1020;
    mem[5681] = 'd1020;
    mem[5682] = 'd1020;
    mem[5683] = 'd1020;
    mem[5684] = 'd1020;
    mem[5685] = 'd1020;
    mem[5686] = 'd1020;
    mem[5687] = 'd1020;
    mem[5688] = 'd1020;
    mem[5689] = 'd1020;
    mem[5690] = 'd1020;
    mem[5691] = 'd1020;
    mem[5692] = 'd1020;
    mem[5693] = 'd1020;
    mem[5694] = 'd1020;
    mem[5695] = 'd1020;
    mem[5696] = 'd1020;
    mem[5697] = 'd1020;
    mem[5698] = 'd1020;
    mem[5699] = 'd1020;
    mem[5700] = 'd1020;
    mem[5701] = 'd1020;
    mem[5702] = 'd1020;
    mem[5703] = 'd1020;
    mem[5704] = 'd1020;
    mem[5705] = 'd1020;
    mem[5706] = 'd1020;
    mem[5707] = 'd1020;
    mem[5708] = 'd1020;
    mem[5709] = 'd1020;
    mem[5710] = 'd1020;
    mem[5711] = 'd1020;
    mem[5712] = 'd1020;
    mem[5713] = 'd1020;
    mem[5714] = 'd1020;
    mem[5715] = 'd1020;
    mem[5716] = 'd1020;
    mem[5717] = 'd1020;
    mem[5718] = 'd1020;
    mem[5719] = 'd1020;
    mem[5720] = 'd1020;
    mem[5721] = 'd1020;
    mem[5722] = 'd1020;
    mem[5723] = 'd1020;
    mem[5724] = 'd1020;
    mem[5725] = 'd1020;
    mem[5726] = 'd1016;
    mem[5727] = 'd1020;
    mem[5728] = 'd1016;
    mem[5729] = 'd1020;
    mem[5730] = 'd1016;
    mem[5731] = 'd1020;
    mem[5732] = 'd1016;
    mem[5733] = 'd1020;
    mem[5734] = 'd1016;
    mem[5735] = 'd1020;
    mem[5736] = 'd1012;
    mem[5737] = 'd1020;
    mem[5738] = 'd1012;
    mem[5739] = 'd1020;
    mem[5740] = 'd1016;
    mem[5741] = 'd1020;
    mem[5742] = 'd1016;
    mem[5743] = 'd1020;
    mem[5744] = 'd1016;
    mem[5745] = 'd1020;
    mem[5746] = 'd1016;
    mem[5747] = 'd1020;
    mem[5748] = 'd1016;
    mem[5749] = 'd1020;
    mem[5750] = 'd1020;
    mem[5751] = 'd1020;
    mem[5752] = 'd1020;
    mem[5753] = 'd1020;
    mem[5754] = 'd1020;
    mem[5755] = 'd1020;
    mem[5756] = 'd1020;
    mem[5757] = 'd1020;
    mem[5758] = 'd1020;
    mem[5759] = 'd1020;
    mem[5760] = 'd1020;
    mem[5761] = 'd1020;
    mem[5762] = 'd1020;
    mem[5763] = 'd1020;
    mem[5764] = 'd1020;
    mem[5765] = 'd1020;
    mem[5766] = 'd1020;
    mem[5767] = 'd1020;
    mem[5768] = 'd1020;
    mem[5769] = 'd1020;
    mem[5770] = 'd1020;
    mem[5771] = 'd1020;
    mem[5772] = 'd1020;
    mem[5773] = 'd1020;
    mem[5774] = 'd1020;
    mem[5775] = 'd1020;

end


endmodule

module image_gen_colorbar #(
    parameter X_RESOLUTION = 1288,
    parameter Y_RESOLUTION = 768,
    parameter H_FRONT_PORCH = 50, // 2x X_RESOLUTION
    parameter H_BACK_PORCH = 50, // ~ 2.2x X_RESOLUTION
    parameter V_FRONT_PORCH = 2,
    parameter V_BACK_PORCH = 2,
    parameter H_SYNC_PULSE_WIDTH = 44,
    parameter V_SYNC_PULSE_WIDTH = 4
) (
    input logic pixel_clock_in,
    input logic reset_n_in,

    output logic [9:0] pixel_data_red_out,
    output logic [9:0] pixel_data_green_out,
    output logic [9:0] pixel_data_blue_out,
    output logic [9:0] pixel_data_out,

    output logic line_valid,
    output logic frame_valid
);

parameter H_START = H_SYNC_PULSE_WIDTH + H_BACK_PORCH;

logic [31:0] x_counter;
logic [31:0] y_counter;
logic [31:0] pixel_counter;

logic [9:0] mem[5927:0];

always @(posedge pixel_clock_in) begin

    if(!reset_n_in) begin

        pixel_data_red_out <= 0;
        pixel_data_green_out <= 0;
        pixel_data_blue_out <= 0;
        line_valid <= 0;
        frame_valid <= 0;

        x_counter <= 0;
        y_counter <= 0;
        pixel_counter <= 0;

    end 

    else begin
            
        // Increment counters
        if (x_counter <= (H_START + X_RESOLUTION + H_FRONT_PORCH)) begin
            x_counter <= x_counter + 1;
        end

        else begin
            x_counter <= 0;

            if (y_counter <= (V_SYNC_PULSE_WIDTH + V_BACK_PORCH + Y_RESOLUTION + V_FRONT_PORCH)) begin
                y_counter <= y_counter + 1;
            end

            else begin
                y_counter <= 0;
            end 

        end

        // Output line valud
        if ((x_counter >= (H_START)) &&
            (x_counter < (H_START + X_RESOLUTION)) &&
            (y_counter >= (V_SYNC_PULSE_WIDTH + V_BACK_PORCH)) &&
            (y_counter < (V_SYNC_PULSE_WIDTH + V_BACK_PORCH + Y_RESOLUTION))) begin
                
            line_valid <= 1;

            pixel_counter <= pixel_counter + 1;

            if ((x_counter >= (H_START)) &&
                (x_counter < (H_START + 100))) begin
                    pixel_data_red_out <= 'h3ff;
                    pixel_data_green_out <= 'h00;
                    pixel_data_blue_out <= 'h00;

                    if (!x_counter[0] && !y_counter[0]) pixel_data_out <= 'h0; //b
                    else if (x_counter[1] && !y_counter[0]) pixel_data_out <= 'h0; //g
                    else if (!x_counter[0] && y_counter[0]) pixel_data_out <= 'h0; //g
                    else if (x_counter[0] && y_counter[0]) pixel_data_out <= 'h3ff; //r
                end
            else if ((x_counter >= (H_START + 100)) &&
                (x_counter < (H_START + 200))) begin
                    pixel_data_red_out <= 'h00;
                    pixel_data_green_out <= 'h3ff;
                    pixel_data_blue_out <= 'h00;

                    if (!x_counter[0] && !y_counter[0]) pixel_data_out <= 'h3ff; //b
                    else if (x_counter[1] && !y_counter[0]) pixel_data_out <= 'h3ff; //g
                    else if (!x_counter[0] && y_counter[0]) pixel_data_out <= 'h3ff; //g
                    else if (x_counter[0] && y_counter[0]) pixel_data_out <= 'h0; //r
                end

            else if ((x_counter >= (H_START + 200)) &&
                (x_counter < (H_START + 300))) begin
                    pixel_data_red_out <= 'h00;
                    pixel_data_green_out <= 'h00;
                    pixel_data_blue_out <= 'h3ff;

                    if (!x_counter[0] && !y_counter[0]) pixel_data_out <= 'h3ff; //b
                    else if (x_counter[1] && !y_counter[0]) pixel_data_out <= 'h0; //g
                    else if (!x_counter[0] && y_counter[0]) pixel_data_out <= 'h0; //g
                    else if (x_counter[0] && y_counter[0]) pixel_data_out <= 'h0; //r
                end

            else if ((x_counter >= (H_START + 300)) &&
                (x_counter < (H_START + 400))) begin
                    pixel_data_red_out <= 'h3ff;
                    pixel_data_green_out <= 'h3ff;
                    pixel_data_blue_out <= 'h00;

                    if (!x_counter[0] && !y_counter[0]) pixel_data_out <= 'h0; //b
                    else if (x_counter[1] && !y_counter[0]) pixel_data_out <= 'h3ff; //g
                    else if (!x_counter[0] && y_counter[0]) pixel_data_out <= 'h3ff; //g
                    else if (x_counter[0] && y_counter[0]) pixel_data_out <= 'h3ff; //r
                end

            else if ((x_counter >= (H_START + 400)) &&
                (x_counter < (H_START + 500))) begin
                    pixel_data_red_out <= 'h00;
                    pixel_data_green_out <= 'h3ff;
                    pixel_data_blue_out <= 'h3ff;

                    if (!x_counter[0] && !y_counter[0]) pixel_data_out <= 'h0; //b
                    else if (x_counter[1] && !y_counter[0]) pixel_data_out <= 'h3ff; //g
                    else if (!x_counter[0] && y_counter[0]) pixel_data_out <= 'h3ff; //g
                    else if (x_counter[0] && y_counter[0]) pixel_data_out <= 'h0; //r
                end

            else if ((x_counter >= (H_START + 500)) &&
                (x_counter < (H_START + 600))) begin
                    pixel_data_red_out <= 'h3ff;
                    pixel_data_green_out <= 'h00;
                    pixel_data_blue_out <= 'h3ff;

                    if (!x_counter[0] && !y_counter[0]) pixel_data_out <= 'h3ff; //b
                    else if (x_counter[1] && !y_counter[0]) pixel_data_out <= 'h0; //g
                    else if (!x_counter[0] && y_counter[0]) pixel_data_out <= 'h0; //g
                    else if (x_counter[0] && y_counter[0]) pixel_data_out <= 'h3ff; //r
                end

            else begin
                    pixel_data_red_out <= 'h3ff;
                    pixel_data_green_out <= 'h3ff;
                    pixel_data_blue_out <= 'h3ff;

                    if (!x_counter[0] && !y_counter[0]) pixel_data_out <= 'h3ff; //b
                    else if (x_counter[1] && !y_counter[0]) pixel_data_out <= 'h3ff; //g
                    else if (!x_counter[0] && y_counter[0]) pixel_data_out <= 'h3ff; //g
                    else if (x_counter[0] && y_counter[0]) pixel_data_out <= 'h3ff; //r
                end

        end

        else begin
            line_valid <= 0;
        end

        // Output frame valid
        if (y_counter >= 0 &&
            y_counter < V_SYNC_PULSE_WIDTH) begin

            frame_valid <= 0;
            pixel_counter <= 0;

        end

        else begin
            frame_valid <= 1;
        end

    end

end

endmodule