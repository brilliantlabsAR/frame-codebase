/*
 * This file is a part of: https://github.com/brilliantlabsAR/frame-codebase
 *
 * Authored by: Rohit Rathnam / Silicon Witchery AB (rohit@siliconwitchery.com)
 *              Raj Nakarja / Brilliant Labs Limited (raj@brilliant.xyz)
 *
 * CERN Open Hardware Licence Version 2 - Permissive
 *
 * Copyright © 2023 Brilliant Labs Limited
 */

`timescale 10ns / 10ns

`include "../graphics.sv"

module graphics_tb;

logic spi_clock = 0;
logic spi_reset_n = 0;
logic display_clock = 0;
logic display_reset_n = 0;

logic [7:0] opcode;
logic opcode_valid = 0;
logic [7:0] operand;
logic operand_valid = 0;
integer operand_count = 0;

localparam  SPI_HALF_PERIOD = 1;

initial begin
    #(20000*SPI_HALF_PERIOD)
    spi_reset_n <= 1;
    display_reset_n <= 1;
    #(10000*SPI_HALF_PERIOD)

    // Clear command
    send_opcode('h10);
    done();
    #(2100000*SPI_HALF_PERIOD)

    // Draw pixels
    send_opcode('h12);
    send_operand('h00); // X pos
    send_operand('h00);
    send_operand('h00); // Y pos
    send_operand('h00);
    send_operand('h00); // Width
    send_operand('d48);
    send_operand('h2); // Total colors
    send_operand('h00); // palette offset
    send_operand('hFF);
    send_operand('hFF);
    send_operand('hFF);
    send_operand('hFF);
    send_operand('hFF);
    send_operand('hFF);
    send_operand('h80);
    send_operand('h00);
    send_operand('h00);
    send_operand('h00);
    send_operand('h00);
    send_operand('h01);
    done();
    #(30000*SPI_HALF_PERIOD)

    // Show command
    send_opcode('h14);
    done();
    #(2000000*SPI_HALF_PERIOD)

    $writememh("simulation/image_buffer.txt", graphics.display_buffers.buffer_b.mem);
    $finish;
end

graphics graphics (
    .spi_clock_in(spi_clock),
    .spi_reset_n_in(spi_reset_n),

    .display_clock_in(display_clock),
    .display_reset_n_in(display_reset_n),

    .op_code_in(opcode),
    .op_code_valid_in(opcode_valid),
    .operand_in(operand),
    .operand_valid_in(operand_valid),
    .operand_count_in(operand_count),

    .display_clock_out(),
    .display_hsync_out(),
    .display_vsync_out(),
    .display_y_out(),
    .display_cb_out(),
    .display_cr_out()
);

initial begin
    forever #SPI_HALF_PERIOD spi_clock <= ~spi_clock;
end

initial begin
    forever #(2*SPI_HALF_PERIOD) display_clock <= ~display_clock;
end

task send_opcode(
    input logic [7:0] data
);
    begin
        opcode <= data;
        opcode_valid <= 1;
        #(64*SPI_HALF_PERIOD);
    end
endtask

task send_operand(
    input logic [7:0] data
);
    begin
        operand <= data;
        operand_valid <= 1;
        operand_count <= operand_count + 1;
        #(64*SPI_HALF_PERIOD);
        operand_valid <= 0;
        #(8*SPI_HALF_PERIOD);
    end
endtask

task done;
    begin
        opcode_valid <= 0;
        operand_valid <= 0;
        operand_count <= 0;
        #(8*SPI_HALF_PERIOD);
    end
endtask

initial begin
    $dumpfile("simulation/graphics_tb.fst");
    $dumpvars(0, graphics_tb);
end

endmodule