initial begin
    $dumpfile("dump.vcd");
    $dumpvars(); 
end
