`ifndef __JLIB_VH__
`define __JLIB_VH__


`define USE_LATTICE_EBR


`endif // __JLIB_VH__
