module huff_tables  (
    input   logic               clk,
    input   logic [7:0]         symbol[1:0],
    input   logic               re[1:0],
    input   logic [1:0]         sel[1:0], //0..DC-Y, 1..DC-UV, 2..AC-Y, 3..AC-UV
    output  logic [4:0]         len[1:0],
    output  logic [15:0]        code[1:0]
);

//0..DC-Y, 1..DC-UV, 2..AC-Y, 3..AC-UV
logic [19:0] ht0[11:0]; /* synthesis syn_romstyle = "Logic" */
logic [19:0] ht1[11:0]; /* synthesis syn_romstyle = "Logic" */
logic [19:0] ht2[255:0]; /* synthesis syn_romstyle = "Logic" */
logic [19:0] ht3[255:0]; /* synthesis syn_romstyle = "Logic" */

logic [19:0] h[1:0];

always_comb  
    for (int i=0; i<2; i++)
        case(sel[i])
        0: h[i] = ht0[symbol[i][3:0]];
        1: h[i] = ht1[symbol[i][3:0]];
        2: h[i] = ht2[symbol[i]];
        3: h[i] = ht3[symbol[i]];
        endcase


always @(posedge clk)  
    for (int i=0; i<2; i++)
        if (re[i]) begin 
            len[i] <= (h[i] >> 16) + 1; // need to add 1 so there is no need to store extra bit
            code[i] <= h[i] & 'hffff;
        end            

always_comb begin
    ht0[4'h 0] = {4'd  1, 12'b 00_0000000000, 4'b0};
    ht0[4'h 1] = {4'd  2, 12'b 010_000000000, 4'b0};
    ht0[4'h 2] = {4'd  2, 12'b 011_000000000, 4'b0};
    ht0[4'h 3] = {4'd  2, 12'b 100_000000000, 4'b0};
    ht0[4'h 4] = {4'd  2, 12'b 101_000000000, 4'b0};
    ht0[4'h 5] = {4'd  2, 12'b 110_000000000, 4'b0};
    ht0[4'h 6] = {4'd  3, 12'b 1110_00000000, 4'b0};
    ht0[4'h 7] = {4'd  4, 12'b 11110_0000000, 4'b0};
    ht0[4'h 8] = {4'd  5, 12'b 111110_000000, 4'b0};
    ht0[4'h 9] = {4'd  6, 12'b 1111110_00000, 4'b0};
    ht0[4'h a] = {4'd  7, 12'b 11111110_0000, 4'b0};
    ht0[4'h b] = {4'd  8, 12'b 111111110_000, 4'b0}; //len=9
end

always_comb begin
    ht1[4'h 0] = {4'd  1, 12'b 00_0000000000, 4'b0};
    ht1[4'h 1] = {4'd  1, 12'b 01_0000000000, 4'b0};
    ht1[4'h 2] = {4'd  1, 12'b 10_0000000000, 4'b0};
    ht1[4'h 3] = {4'd  2, 12'b 110_000000000, 4'b0};
    ht1[4'h 4] = {4'd  3, 12'b 1110_00000000, 4'b0};
    ht1[4'h 5] = {4'd  4, 12'b 11110_0000000, 4'b0};
    ht1[4'h 6] = {4'd  5, 12'b 111110_000000, 4'b0};
    ht1[4'h 7] = {4'd  6, 12'b 1111110_00000, 4'b0};
    ht1[4'h 8] = {4'd  7, 12'b 11111110_0000, 4'b0};
    ht1[4'h 9] = {4'd  8, 12'b 111111110_000, 4'b0};
    ht1[4'h a] = {4'd  9, 12'b 1111111110_00, 4'b0};
    ht1[4'h b] = {4'd 10, 12'b 11111111110_0, 4'b0}; //len=11
end

always_comb begin
    for (int i=0; i<256; i++) ht2[i] =  20'h x;
    ht2[8'h 01] = {4'd  1, 16'b 00_00000000000000};
    ht2[8'h 02] = {4'd  1, 16'b 01_00000000000000};
    ht2[8'h 03] = {4'd  2, 16'b 100_0000000000000};
    ht2[8'h 00] = {4'd  3, 16'b 1010_000000000000};
    ht2[8'h 04] = {4'd  3, 16'b 1011_000000000000};
    ht2[8'h 11] = {4'd  3, 16'b 1100_000000000000};
    ht2[8'h 05] = {4'd  4, 16'b 11010_00000000000};
    ht2[8'h 12] = {4'd  4, 16'b 11011_00000000000};
    ht2[8'h 21] = {4'd  4, 16'b 11100_00000000000};
    ht2[8'h 31] = {4'd  5, 16'b 111010_0000000000};
    ht2[8'h 41] = {4'd  5, 16'b 111011_0000000000};
    ht2[8'h 06] = {4'd  6, 16'b 1111000_000000000};
    ht2[8'h 13] = {4'd  6, 16'b 1111001_000000000};
    ht2[8'h 51] = {4'd  6, 16'b 1111010_000000000};
    ht2[8'h 61] = {4'd  6, 16'b 1111011_000000000};
    ht2[8'h 07] = {4'd  7, 16'b 11111000_00000000};
    ht2[8'h 22] = {4'd  7, 16'b 11111001_00000000};
    ht2[8'h 71] = {4'd  7, 16'b 11111010_00000000};
    ht2[8'h 14] = {4'd  8, 16'b 111110110_0000000};
    ht2[8'h 32] = {4'd  8, 16'b 111110111_0000000};
    ht2[8'h 81] = {4'd  8, 16'b 111111000_0000000};
    ht2[8'h 91] = {4'd  8, 16'b 111111001_0000000};
    ht2[8'h a1] = {4'd  8, 16'b 111111010_0000000};
    ht2[8'h 08] = {4'd  9, 16'b 1111110110_000000};
    ht2[8'h 23] = {4'd  9, 16'b 1111110111_000000};
    ht2[8'h 42] = {4'd  9, 16'b 1111111000_000000};
    ht2[8'h b1] = {4'd  9, 16'b 1111111001_000000};
    ht2[8'h c1] = {4'd  9, 16'b 1111111010_000000};
    ht2[8'h 15] = {4'd 10, 16'b 11111110110_00000};
    ht2[8'h 52] = {4'd 10, 16'b 11111110111_00000};
    ht2[8'h d1] = {4'd 10, 16'b 11111111000_00000};
    ht2[8'h f0] = {4'd 10, 16'b 11111111001_00000};
    ht2[8'h 24] = {4'd 11, 16'b 111111110100_0000};
    ht2[8'h 33] = {4'd 11, 16'b 111111110101_0000};
    ht2[8'h 62] = {4'd 11, 16'b 111111110110_0000};
    ht2[8'h 72] = {4'd 11, 16'b 111111110111_0000};
    ht2[8'h 82] = {4'd 14, 16'b 111111111000000_0};
    ht2[8'h 09] = {4'd 15, 16'b 1111111110000010};
    ht2[8'h 0a] = {4'd 15, 16'b 1111111110000011};
    ht2[8'h 16] = {4'd 15, 16'b 1111111110000100};
    ht2[8'h 17] = {4'd 15, 16'b 1111111110000101};
    ht2[8'h 18] = {4'd 15, 16'b 1111111110000110};
    ht2[8'h 19] = {4'd 15, 16'b 1111111110000111};
    ht2[8'h 1a] = {4'd 15, 16'b 1111111110001000};
    ht2[8'h 25] = {4'd 15, 16'b 1111111110001001};
    ht2[8'h 26] = {4'd 15, 16'b 1111111110001010};
    ht2[8'h 27] = {4'd 15, 16'b 1111111110001011};
    ht2[8'h 28] = {4'd 15, 16'b 1111111110001100};
    ht2[8'h 29] = {4'd 15, 16'b 1111111110001101};
    ht2[8'h 2a] = {4'd 15, 16'b 1111111110001110};
    ht2[8'h 34] = {4'd 15, 16'b 1111111110001111};
    ht2[8'h 35] = {4'd 15, 16'b 1111111110010000};
    ht2[8'h 36] = {4'd 15, 16'b 1111111110010001};
    ht2[8'h 37] = {4'd 15, 16'b 1111111110010010};
    ht2[8'h 38] = {4'd 15, 16'b 1111111110010011};
    ht2[8'h 39] = {4'd 15, 16'b 1111111110010100};
    ht2[8'h 3a] = {4'd 15, 16'b 1111111110010101};
    ht2[8'h 43] = {4'd 15, 16'b 1111111110010110};
    ht2[8'h 44] = {4'd 15, 16'b 1111111110010111};
    ht2[8'h 45] = {4'd 15, 16'b 1111111110011000};
    ht2[8'h 46] = {4'd 15, 16'b 1111111110011001};
    ht2[8'h 47] = {4'd 15, 16'b 1111111110011010};
    ht2[8'h 48] = {4'd 15, 16'b 1111111110011011};
    ht2[8'h 49] = {4'd 15, 16'b 1111111110011100};
    ht2[8'h 4a] = {4'd 15, 16'b 1111111110011101};
    ht2[8'h 53] = {4'd 15, 16'b 1111111110011110};
    ht2[8'h 54] = {4'd 15, 16'b 1111111110011111};
    ht2[8'h 55] = {4'd 15, 16'b 1111111110100000};
    ht2[8'h 56] = {4'd 15, 16'b 1111111110100001};
    ht2[8'h 57] = {4'd 15, 16'b 1111111110100010};
    ht2[8'h 58] = {4'd 15, 16'b 1111111110100011};
    ht2[8'h 59] = {4'd 15, 16'b 1111111110100100};
    ht2[8'h 5a] = {4'd 15, 16'b 1111111110100101};
    ht2[8'h 63] = {4'd 15, 16'b 1111111110100110};
    ht2[8'h 64] = {4'd 15, 16'b 1111111110100111};
    ht2[8'h 65] = {4'd 15, 16'b 1111111110101000};
    ht2[8'h 66] = {4'd 15, 16'b 1111111110101001};
    ht2[8'h 67] = {4'd 15, 16'b 1111111110101010};
    ht2[8'h 68] = {4'd 15, 16'b 1111111110101011};
    ht2[8'h 69] = {4'd 15, 16'b 1111111110101100};
    ht2[8'h 6a] = {4'd 15, 16'b 1111111110101101};
    ht2[8'h 73] = {4'd 15, 16'b 1111111110101110};
    ht2[8'h 74] = {4'd 15, 16'b 1111111110101111};
    ht2[8'h 75] = {4'd 15, 16'b 1111111110110000};
    ht2[8'h 76] = {4'd 15, 16'b 1111111110110001};
    ht2[8'h 77] = {4'd 15, 16'b 1111111110110010};
    ht2[8'h 78] = {4'd 15, 16'b 1111111110110011};
    ht2[8'h 79] = {4'd 15, 16'b 1111111110110100};
    ht2[8'h 7a] = {4'd 15, 16'b 1111111110110101};
    ht2[8'h 83] = {4'd 15, 16'b 1111111110110110};
    ht2[8'h 84] = {4'd 15, 16'b 1111111110110111};
    ht2[8'h 85] = {4'd 15, 16'b 1111111110111000};
    ht2[8'h 86] = {4'd 15, 16'b 1111111110111001};
    ht2[8'h 87] = {4'd 15, 16'b 1111111110111010};
    ht2[8'h 88] = {4'd 15, 16'b 1111111110111011};
    ht2[8'h 89] = {4'd 15, 16'b 1111111110111100};
    ht2[8'h 8a] = {4'd 15, 16'b 1111111110111101};
    ht2[8'h 92] = {4'd 15, 16'b 1111111110111110};
    ht2[8'h 93] = {4'd 15, 16'b 1111111110111111};
    ht2[8'h 94] = {4'd 15, 16'b 1111111111000000};
    ht2[8'h 95] = {4'd 15, 16'b 1111111111000001};
    ht2[8'h 96] = {4'd 15, 16'b 1111111111000010};
    ht2[8'h 97] = {4'd 15, 16'b 1111111111000011};
    ht2[8'h 98] = {4'd 15, 16'b 1111111111000100};
    ht2[8'h 99] = {4'd 15, 16'b 1111111111000101};
    ht2[8'h 9a] = {4'd 15, 16'b 1111111111000110};
    ht2[8'h a2] = {4'd 15, 16'b 1111111111000111};
    ht2[8'h a3] = {4'd 15, 16'b 1111111111001000};
    ht2[8'h a4] = {4'd 15, 16'b 1111111111001001};
    ht2[8'h a5] = {4'd 15, 16'b 1111111111001010};
    ht2[8'h a6] = {4'd 15, 16'b 1111111111001011};
    ht2[8'h a7] = {4'd 15, 16'b 1111111111001100};
    ht2[8'h a8] = {4'd 15, 16'b 1111111111001101};
    ht2[8'h a9] = {4'd 15, 16'b 1111111111001110};
    ht2[8'h aa] = {4'd 15, 16'b 1111111111001111};
    ht2[8'h b2] = {4'd 15, 16'b 1111111111010000};
    ht2[8'h b3] = {4'd 15, 16'b 1111111111010001};
    ht2[8'h b4] = {4'd 15, 16'b 1111111111010010};
    ht2[8'h b5] = {4'd 15, 16'b 1111111111010011};
    ht2[8'h b6] = {4'd 15, 16'b 1111111111010100};
    ht2[8'h b7] = {4'd 15, 16'b 1111111111010101};
    ht2[8'h b8] = {4'd 15, 16'b 1111111111010110};
    ht2[8'h b9] = {4'd 15, 16'b 1111111111010111};
    ht2[8'h ba] = {4'd 15, 16'b 1111111111011000};
    ht2[8'h c2] = {4'd 15, 16'b 1111111111011001};
    ht2[8'h c3] = {4'd 15, 16'b 1111111111011010};
    ht2[8'h c4] = {4'd 15, 16'b 1111111111011011};
    ht2[8'h c5] = {4'd 15, 16'b 1111111111011100};
    ht2[8'h c6] = {4'd 15, 16'b 1111111111011101};
    ht2[8'h c7] = {4'd 15, 16'b 1111111111011110};
    ht2[8'h c8] = {4'd 15, 16'b 1111111111011111};
    ht2[8'h c9] = {4'd 15, 16'b 1111111111100000};
    ht2[8'h ca] = {4'd 15, 16'b 1111111111100001};
    ht2[8'h d2] = {4'd 15, 16'b 1111111111100010};
    ht2[8'h d3] = {4'd 15, 16'b 1111111111100011};
    ht2[8'h d4] = {4'd 15, 16'b 1111111111100100};
    ht2[8'h d5] = {4'd 15, 16'b 1111111111100101};
    ht2[8'h d6] = {4'd 15, 16'b 1111111111100110};
    ht2[8'h d7] = {4'd 15, 16'b 1111111111100111};
    ht2[8'h d8] = {4'd 15, 16'b 1111111111101000};
    ht2[8'h d9] = {4'd 15, 16'b 1111111111101001};
    ht2[8'h da] = {4'd 15, 16'b 1111111111101010};
    ht2[8'h e1] = {4'd 15, 16'b 1111111111101011};
    ht2[8'h e2] = {4'd 15, 16'b 1111111111101100};
    ht2[8'h e3] = {4'd 15, 16'b 1111111111101101};
    ht2[8'h e4] = {4'd 15, 16'b 1111111111101110};
    ht2[8'h e5] = {4'd 15, 16'b 1111111111101111};
    ht2[8'h e6] = {4'd 15, 16'b 1111111111110000};
    ht2[8'h e7] = {4'd 15, 16'b 1111111111110001};
    ht2[8'h e8] = {4'd 15, 16'b 1111111111110010};
    ht2[8'h e9] = {4'd 15, 16'b 1111111111110011};
    ht2[8'h ea] = {4'd 15, 16'b 1111111111110100};
    ht2[8'h f1] = {4'd 15, 16'b 1111111111110101};
    ht2[8'h f2] = {4'd 15, 16'b 1111111111110110};
    ht2[8'h f3] = {4'd 15, 16'b 1111111111110111};
    ht2[8'h f4] = {4'd 15, 16'b 1111111111111000};
    ht2[8'h f5] = {4'd 15, 16'b 1111111111111001};
    ht2[8'h f6] = {4'd 15, 16'b 1111111111111010};
    ht2[8'h f7] = {4'd 15, 16'b 1111111111111011};
    ht2[8'h f8] = {4'd 15, 16'b 1111111111111100};
    ht2[8'h f9] = {4'd 15, 16'b 1111111111111101};
    ht2[8'h fa] = {4'd 15, 16'b 1111111111111110};
end

always_comb begin
    for (int i=0; i<256; i++) ht3[i] =  20'h x;
    ht3[8'h 00] = {4'd  1, 16'b 00_00000000000000};
    ht3[8'h 01] = {4'd  1, 16'b 01_00000000000000};
    ht3[8'h 02] = {4'd  2, 16'b 100_0000000000000};
    ht3[8'h 03] = {4'd  3, 16'b 1010_000000000000};
    ht3[8'h 11] = {4'd  3, 16'b 1011_000000000000};
    ht3[8'h 04] = {4'd  4, 16'b 11000_00000000000};
    ht3[8'h 05] = {4'd  4, 16'b 11001_00000000000};
    ht3[8'h 21] = {4'd  4, 16'b 11010_00000000000};
    ht3[8'h 31] = {4'd  4, 16'b 11011_00000000000};
    ht3[8'h 06] = {4'd  5, 16'b 111000_0000000000};
    ht3[8'h 12] = {4'd  5, 16'b 111001_0000000000};
    ht3[8'h 41] = {4'd  5, 16'b 111010_0000000000};
    ht3[8'h 51] = {4'd  5, 16'b 111011_0000000000};
    ht3[8'h 07] = {4'd  6, 16'b 1111000_000000000};
    ht3[8'h 61] = {4'd  6, 16'b 1111001_000000000};
    ht3[8'h 71] = {4'd  6, 16'b 1111010_000000000};
    ht3[8'h 13] = {4'd  7, 16'b 11110110_00000000};
    ht3[8'h 22] = {4'd  7, 16'b 11110111_00000000};
    ht3[8'h 32] = {4'd  7, 16'b 11111000_00000000};
    ht3[8'h 81] = {4'd  7, 16'b 11111001_00000000};
    ht3[8'h 08] = {4'd  8, 16'b 111110100_0000000};
    ht3[8'h 14] = {4'd  8, 16'b 111110101_0000000};
    ht3[8'h 42] = {4'd  8, 16'b 111110110_0000000};
    ht3[8'h 91] = {4'd  8, 16'b 111110111_0000000};
    ht3[8'h a1] = {4'd  8, 16'b 111111000_0000000};
    ht3[8'h b1] = {4'd  8, 16'b 111111001_0000000};
    ht3[8'h c1] = {4'd  8, 16'b 111111010_0000000};
    ht3[8'h 09] = {4'd  9, 16'b 1111110110_000000};
    ht3[8'h 23] = {4'd  9, 16'b 1111110111_000000};
    ht3[8'h 33] = {4'd  9, 16'b 1111111000_000000};
    ht3[8'h 52] = {4'd  9, 16'b 1111111001_000000};
    ht3[8'h f0] = {4'd  9, 16'b 1111111010_000000};
    ht3[8'h 15] = {4'd 10, 16'b 11111110110_00000};
    ht3[8'h 62] = {4'd 10, 16'b 11111110111_00000};
    ht3[8'h 72] = {4'd 10, 16'b 11111111000_00000};
    ht3[8'h d1] = {4'd 10, 16'b 11111111001_00000};
    ht3[8'h 0a] = {4'd 11, 16'b 111111110100_0000};
    ht3[8'h 16] = {4'd 11, 16'b 111111110101_0000};
    ht3[8'h 24] = {4'd 11, 16'b 111111110110_0000};
    ht3[8'h 34] = {4'd 11, 16'b 111111110111_0000};
    ht3[8'h e1] = {4'd 13, 16'b 11111111100000_00};
    ht3[8'h 25] = {4'd 14, 16'b 111111111000010_0};
    ht3[8'h f1] = {4'd 14, 16'b 111111111000011_0};
    ht3[8'h 17] = {4'd 15, 16'b 1111111110001000};
    ht3[8'h 18] = {4'd 15, 16'b 1111111110001001};
    ht3[8'h 19] = {4'd 15, 16'b 1111111110001010};
    ht3[8'h 1a] = {4'd 15, 16'b 1111111110001011};
    ht3[8'h 26] = {4'd 15, 16'b 1111111110001100};
    ht3[8'h 27] = {4'd 15, 16'b 1111111110001101};
    ht3[8'h 28] = {4'd 15, 16'b 1111111110001110};
    ht3[8'h 29] = {4'd 15, 16'b 1111111110001111};
    ht3[8'h 2a] = {4'd 15, 16'b 1111111110010000};
    ht3[8'h 35] = {4'd 15, 16'b 1111111110010001};
    ht3[8'h 36] = {4'd 15, 16'b 1111111110010010};
    ht3[8'h 37] = {4'd 15, 16'b 1111111110010011};
    ht3[8'h 38] = {4'd 15, 16'b 1111111110010100};
    ht3[8'h 39] = {4'd 15, 16'b 1111111110010101};
    ht3[8'h 3a] = {4'd 15, 16'b 1111111110010110};
    ht3[8'h 43] = {4'd 15, 16'b 1111111110010111};
    ht3[8'h 44] = {4'd 15, 16'b 1111111110011000};
    ht3[8'h 45] = {4'd 15, 16'b 1111111110011001};
    ht3[8'h 46] = {4'd 15, 16'b 1111111110011010};
    ht3[8'h 47] = {4'd 15, 16'b 1111111110011011};
    ht3[8'h 48] = {4'd 15, 16'b 1111111110011100};
    ht3[8'h 49] = {4'd 15, 16'b 1111111110011101};
    ht3[8'h 4a] = {4'd 15, 16'b 1111111110011110};
    ht3[8'h 53] = {4'd 15, 16'b 1111111110011111};
    ht3[8'h 54] = {4'd 15, 16'b 1111111110100000};
    ht3[8'h 55] = {4'd 15, 16'b 1111111110100001};
    ht3[8'h 56] = {4'd 15, 16'b 1111111110100010};
    ht3[8'h 57] = {4'd 15, 16'b 1111111110100011};
    ht3[8'h 58] = {4'd 15, 16'b 1111111110100100};
    ht3[8'h 59] = {4'd 15, 16'b 1111111110100101};
    ht3[8'h 5a] = {4'd 15, 16'b 1111111110100110};
    ht3[8'h 63] = {4'd 15, 16'b 1111111110100111};
    ht3[8'h 64] = {4'd 15, 16'b 1111111110101000};
    ht3[8'h 65] = {4'd 15, 16'b 1111111110101001};
    ht3[8'h 66] = {4'd 15, 16'b 1111111110101010};
    ht3[8'h 67] = {4'd 15, 16'b 1111111110101011};
    ht3[8'h 68] = {4'd 15, 16'b 1111111110101100};
    ht3[8'h 69] = {4'd 15, 16'b 1111111110101101};
    ht3[8'h 6a] = {4'd 15, 16'b 1111111110101110};
    ht3[8'h 73] = {4'd 15, 16'b 1111111110101111};
    ht3[8'h 74] = {4'd 15, 16'b 1111111110110000};
    ht3[8'h 75] = {4'd 15, 16'b 1111111110110001};
    ht3[8'h 76] = {4'd 15, 16'b 1111111110110010};
    ht3[8'h 77] = {4'd 15, 16'b 1111111110110011};
    ht3[8'h 78] = {4'd 15, 16'b 1111111110110100};
    ht3[8'h 79] = {4'd 15, 16'b 1111111110110101};
    ht3[8'h 7a] = {4'd 15, 16'b 1111111110110110};
    ht3[8'h 82] = {4'd 15, 16'b 1111111110110111};
    ht3[8'h 83] = {4'd 15, 16'b 1111111110111000};
    ht3[8'h 84] = {4'd 15, 16'b 1111111110111001};
    ht3[8'h 85] = {4'd 15, 16'b 1111111110111010};
    ht3[8'h 86] = {4'd 15, 16'b 1111111110111011};
    ht3[8'h 87] = {4'd 15, 16'b 1111111110111100};
    ht3[8'h 88] = {4'd 15, 16'b 1111111110111101};
    ht3[8'h 89] = {4'd 15, 16'b 1111111110111110};
    ht3[8'h 8a] = {4'd 15, 16'b 1111111110111111};
    ht3[8'h 92] = {4'd 15, 16'b 1111111111000000};
    ht3[8'h 93] = {4'd 15, 16'b 1111111111000001};
    ht3[8'h 94] = {4'd 15, 16'b 1111111111000010};
    ht3[8'h 95] = {4'd 15, 16'b 1111111111000011};
    ht3[8'h 96] = {4'd 15, 16'b 1111111111000100};
    ht3[8'h 97] = {4'd 15, 16'b 1111111111000101};
    ht3[8'h 98] = {4'd 15, 16'b 1111111111000110};
    ht3[8'h 99] = {4'd 15, 16'b 1111111111000111};
    ht3[8'h 9a] = {4'd 15, 16'b 1111111111001000};
    ht3[8'h a2] = {4'd 15, 16'b 1111111111001001};
    ht3[8'h a3] = {4'd 15, 16'b 1111111111001010};
    ht3[8'h a4] = {4'd 15, 16'b 1111111111001011};
    ht3[8'h a5] = {4'd 15, 16'b 1111111111001100};
    ht3[8'h a6] = {4'd 15, 16'b 1111111111001101};
    ht3[8'h a7] = {4'd 15, 16'b 1111111111001110};
    ht3[8'h a8] = {4'd 15, 16'b 1111111111001111};
    ht3[8'h a9] = {4'd 15, 16'b 1111111111010000};
    ht3[8'h aa] = {4'd 15, 16'b 1111111111010001};
    ht3[8'h b2] = {4'd 15, 16'b 1111111111010010};
    ht3[8'h b3] = {4'd 15, 16'b 1111111111010011};
    ht3[8'h b4] = {4'd 15, 16'b 1111111111010100};
    ht3[8'h b5] = {4'd 15, 16'b 1111111111010101};
    ht3[8'h b6] = {4'd 15, 16'b 1111111111010110};
    ht3[8'h b7] = {4'd 15, 16'b 1111111111010111};
    ht3[8'h b8] = {4'd 15, 16'b 1111111111011000};
    ht3[8'h b9] = {4'd 15, 16'b 1111111111011001};
    ht3[8'h ba] = {4'd 15, 16'b 1111111111011010};
    ht3[8'h c2] = {4'd 15, 16'b 1111111111011011};
    ht3[8'h c3] = {4'd 15, 16'b 1111111111011100};
    ht3[8'h c4] = {4'd 15, 16'b 1111111111011101};
    ht3[8'h c5] = {4'd 15, 16'b 1111111111011110};
    ht3[8'h c6] = {4'd 15, 16'b 1111111111011111};
    ht3[8'h c7] = {4'd 15, 16'b 1111111111100000};
    ht3[8'h c8] = {4'd 15, 16'b 1111111111100001};
    ht3[8'h c9] = {4'd 15, 16'b 1111111111100010};
    ht3[8'h ca] = {4'd 15, 16'b 1111111111100011};
    ht3[8'h d2] = {4'd 15, 16'b 1111111111100100};
    ht3[8'h d3] = {4'd 15, 16'b 1111111111100101};
    ht3[8'h d4] = {4'd 15, 16'b 1111111111100110};
    ht3[8'h d5] = {4'd 15, 16'b 1111111111100111};
    ht3[8'h d6] = {4'd 15, 16'b 1111111111101000};
    ht3[8'h d7] = {4'd 15, 16'b 1111111111101001};
    ht3[8'h d8] = {4'd 15, 16'b 1111111111101010};
    ht3[8'h d9] = {4'd 15, 16'b 1111111111101011};
    ht3[8'h da] = {4'd 15, 16'b 1111111111101100};
    ht3[8'h e2] = {4'd 15, 16'b 1111111111101101};
    ht3[8'h e3] = {4'd 15, 16'b 1111111111101110};
    ht3[8'h e4] = {4'd 15, 16'b 1111111111101111};
    ht3[8'h e5] = {4'd 15, 16'b 1111111111110000};
    ht3[8'h e6] = {4'd 15, 16'b 1111111111110001};
    ht3[8'h e7] = {4'd 15, 16'b 1111111111110010};
    ht3[8'h e8] = {4'd 15, 16'b 1111111111110011};
    ht3[8'h e9] = {4'd 15, 16'b 1111111111110100};
    ht3[8'h ea] = {4'd 15, 16'b 1111111111110101};
    ht3[8'h f2] = {4'd 15, 16'b 1111111111110110};
    ht3[8'h f3] = {4'd 15, 16'b 1111111111110111};
    ht3[8'h f4] = {4'd 15, 16'b 1111111111111000};
    ht3[8'h f5] = {4'd 15, 16'b 1111111111111001};
    ht3[8'h f6] = {4'd 15, 16'b 1111111111111010};
    ht3[8'h f7] = {4'd 15, 16'b 1111111111111011};
    ht3[8'h f8] = {4'd 15, 16'b 1111111111111100};
    ht3[8'h f9] = {4'd 15, 16'b 1111111111111101};
    ht3[8'h fa] = {4'd 15, 16'b 1111111111111110};
end
endmodule
