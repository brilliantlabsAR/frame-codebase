/*
 * This file is a part of: https://github.com/brilliantlabsAR/frame-codebase
 *
 * Authored by: Rohit Rathnam / Silicon Witchery AB (rohit@siliconwitchery.com)
 *              Raj Nakarja / Brilliant Labs Limited (raj@brilliant.xyz)
 *
 * CERN Open Hardware Licence Version 2 - Permissive
 *
 * Copyright © 2023 Brilliant Labs Limited
 */

module image_gen #(
    parameter X_RESOLUTION = 78,
    parameter Y_RESOLUTION = 76,
    parameter H_FRONT_PORCH = 156, // 2x X_RESOLUTION
    parameter H_BACK_PORCH = 172, // ~ 2.2x X_RESOLUTION
    parameter V_FRONT_PORCH = 1,
    parameter V_BACK_PORCH = 2,
    parameter H_SYNC_PULSE_WIDTH = 44,
    parameter V_SYNC_PULSE_WIDTH = 5
) (
    input logic pixel_clock_in,
    input logic reset_n_in,

    output logic [9:0] pixel_data_out,
    output logic line_valid,
    output logic frame_valid
);

logic [31:0] x_counter;
logic [31:0] y_counter;
logic [31:0] pixel_counter;

logic [9:0] mem[17783:0];

always @(posedge pixel_clock_in) begin

    if(!reset_n_in) begin

        pixel_data_out <= 0;
        line_valid <= 0;
        frame_valid <= 0;

        x_counter <= 0;
        y_counter <= 0;
        pixel_counter <= 0;

    end 

    else begin
            
        // Increment counters
        if (x_counter <= (H_SYNC_PULSE_WIDTH + H_BACK_PORCH + X_RESOLUTION + H_FRONT_PORCH)) begin
            x_counter <= x_counter + 1;
        end

        else begin
            x_counter <= 0;

            if (y_counter <= (V_SYNC_PULSE_WIDTH + V_BACK_PORCH + Y_RESOLUTION + V_FRONT_PORCH)) begin
                y_counter <= y_counter + 1;
            end

            else begin
                y_counter <= 0;
            end 

        end

        // Output line valud
        if ((x_counter >= (H_SYNC_PULSE_WIDTH + H_BACK_PORCH)) &&
            (x_counter < (H_SYNC_PULSE_WIDTH + H_BACK_PORCH + X_RESOLUTION)) &&
            (y_counter >= (V_SYNC_PULSE_WIDTH + V_BACK_PORCH)) &&
            (y_counter < (V_SYNC_PULSE_WIDTH + V_BACK_PORCH + Y_RESOLUTION))) begin
                
            line_valid <= 1;

            pixel_counter <= pixel_counter + 1;
        end

        else begin
            line_valid <= 0;
        end

        // Output frame valid
        if (y_counter >= 0 &&
            y_counter < V_SYNC_PULSE_WIDTH) begin

            frame_valid <= 0;
            pixel_counter <= 0;

        end

        else begin
            frame_valid <= 1;
        end
        
        // Output pixel
        pixel_data_out <= mem[pixel_counter];

    end

end

initial begin

    mem[0] = 'd0;
    mem[1] = 'd0;
    mem[2] = 'd1020;
    mem[3] = 'd0;
    mem[4] = 'd1020;
    mem[5] = 'd0;
    mem[6] = 'd0;
    mem[7] = 'd0;
    mem[8] = 'd1020;
    mem[9] = 'd0;
    mem[10] = 'd1020;
    mem[11] = 'd0;
    mem[12] = 'd0;
    mem[13] = 'd0;
    mem[14] = 'd1020;
    mem[15] = 'd0;
    mem[16] = 'd1020;
    mem[17] = 'd0;
    mem[18] = 'd0;
    mem[19] = 'd0;
    mem[20] = 'd1020;
    mem[21] = 'd0;
    mem[22] = 'd1020;
    mem[23] = 'd0;
    mem[24] = 'd0;
    mem[25] = 'd0;
    mem[26] = 'd1020;
    mem[27] = 'd0;
    mem[28] = 'd1020;
    mem[29] = 'd0;
    mem[30] = 'd0;
    mem[31] = 'd0;
    mem[32] = 'd1020;
    mem[33] = 'd0;
    mem[34] = 'd1020;
    mem[35] = 'd0;
    mem[36] = 'd0;
    mem[37] = 'd0;
    mem[38] = 'd1020;
    mem[39] = 'd0;
    mem[40] = 'd1020;
    mem[41] = 'd0;
    mem[42] = 'd0;
    mem[43] = 'd0;
    mem[44] = 'd1020;
    mem[45] = 'd0;
    mem[46] = 'd1020;
    mem[47] = 'd0;
    mem[48] = 'd0;
    mem[49] = 'd0;
    mem[50] = 'd1020;
    mem[51] = 'd0;
    mem[52] = 'd1020;
    mem[53] = 'd0;
    mem[54] = 'd0;
    mem[55] = 'd0;
    mem[56] = 'd1020;
    mem[57] = 'd0;
    mem[58] = 'd1020;
    mem[59] = 'd0;
    mem[60] = 'd0;
    mem[61] = 'd0;
    mem[62] = 'd1020;
    mem[63] = 'd0;
    mem[64] = 'd1020;
    mem[65] = 'd0;
    mem[66] = 'd0;
    mem[67] = 'd0;
    mem[68] = 'd1020;
    mem[69] = 'd0;
    mem[70] = 'd1020;
    mem[71] = 'd0;
    mem[72] = 'd0;
    mem[73] = 'd0;
    mem[74] = 'd1020;
    mem[75] = 'd0;
    mem[76] = 'd1020;
    mem[77] = 'd0;
    mem[78] = 'd0;
    mem[79] = 'd0;
    mem[80] = 'd1020;
    mem[81] = 'd0;
    mem[82] = 'd1020;
    mem[83] = 'd0;
    mem[84] = 'd0;
    mem[85] = 'd0;
    mem[86] = 'd1020;
    mem[87] = 'd0;
    mem[88] = 'd1020;
    mem[89] = 'd0;
    mem[90] = 'd0;
    mem[91] = 'd0;
    mem[92] = 'd1020;
    mem[93] = 'd0;
    mem[94] = 'd1020;
    mem[95] = 'd0;
    mem[96] = 'd0;
    mem[97] = 'd0;
    mem[98] = 'd1020;
    mem[99] = 'd0;
    mem[100] = 'd1020;
    mem[101] = 'd0;
    mem[102] = 'd0;
    mem[103] = 'd0;
    mem[104] = 'd1020;
    mem[105] = 'd0;
    mem[106] = 'd1020;
    mem[107] = 'd0;
    mem[108] = 'd0;
    mem[109] = 'd0;
    mem[110] = 'd1020;
    mem[111] = 'd0;
    mem[112] = 'd1020;
    mem[113] = 'd0;
    mem[114] = 'd0;
    mem[115] = 'd0;
    mem[116] = 'd1020;
    mem[117] = 'd0;
    mem[118] = 'd1020;
    mem[119] = 'd0;
    mem[120] = 'd0;
    mem[121] = 'd0;
    mem[122] = 'd1020;
    mem[123] = 'd0;
    mem[124] = 'd1020;
    mem[125] = 'd0;
    mem[126] = 'd0;
    mem[127] = 'd0;
    mem[128] = 'd1020;
    mem[129] = 'd0;
    mem[130] = 'd1020;
    mem[131] = 'd0;
    mem[132] = 'd0;
    mem[133] = 'd0;
    mem[134] = 'd1020;
    mem[135] = 'd0;
    mem[136] = 'd1020;
    mem[137] = 'd0;
    mem[138] = 'd0;
    mem[139] = 'd0;
    mem[140] = 'd1020;
    mem[141] = 'd0;
    mem[142] = 'd1020;
    mem[143] = 'd0;
    mem[144] = 'd0;
    mem[145] = 'd0;
    mem[146] = 'd1020;
    mem[147] = 'd0;
    mem[148] = 'd1020;
    mem[149] = 'd0;
    mem[150] = 'd0;
    mem[151] = 'd0;
    mem[152] = 'd1020;
    mem[153] = 'd0;
    mem[154] = 'd1020;
    mem[155] = 'd0;
    mem[156] = 'd0;
    mem[157] = 'd0;
    mem[158] = 'd1020;
    mem[159] = 'd0;
    mem[160] = 'd1020;
    mem[161] = 'd0;
    mem[162] = 'd0;
    mem[163] = 'd0;
    mem[164] = 'd1020;
    mem[165] = 'd0;
    mem[166] = 'd1020;
    mem[167] = 'd0;
    mem[168] = 'd0;
    mem[169] = 'd0;
    mem[170] = 'd1020;
    mem[171] = 'd0;
    mem[172] = 'd1020;
    mem[173] = 'd0;
    mem[174] = 'd0;
    mem[175] = 'd0;
    mem[176] = 'd1020;
    mem[177] = 'd0;
    mem[178] = 'd1020;
    mem[179] = 'd0;
    mem[180] = 'd0;
    mem[181] = 'd0;
    mem[182] = 'd1020;
    mem[183] = 'd0;
    mem[184] = 'd1020;
    mem[185] = 'd0;
    mem[186] = 'd0;
    mem[187] = 'd0;
    mem[188] = 'd1020;
    mem[189] = 'd0;
    mem[190] = 'd1020;
    mem[191] = 'd0;
    mem[192] = 'd0;
    mem[193] = 'd0;
    mem[194] = 'd1020;
    mem[195] = 'd0;
    mem[196] = 'd1020;
    mem[197] = 'd0;
    mem[198] = 'd0;
    mem[199] = 'd0;
    mem[200] = 'd1020;
    mem[201] = 'd0;
    mem[202] = 'd1020;
    mem[203] = 'd0;
    mem[204] = 'd0;
    mem[205] = 'd0;
    mem[206] = 'd1020;
    mem[207] = 'd0;
    mem[208] = 'd1020;
    mem[209] = 'd0;
    mem[210] = 'd0;
    mem[211] = 'd0;
    mem[212] = 'd1020;
    mem[213] = 'd0;
    mem[214] = 'd1020;
    mem[215] = 'd0;
    mem[216] = 'd0;
    mem[217] = 'd0;
    mem[218] = 'd1020;
    mem[219] = 'd0;
    mem[220] = 'd1020;
    mem[221] = 'd0;
    mem[222] = 'd0;
    mem[223] = 'd0;
    mem[224] = 'd1020;
    mem[225] = 'd0;
    mem[226] = 'd1020;
    mem[227] = 'd0;
    mem[228] = 'd0;
    mem[229] = 'd0;
    mem[230] = 'd1020;
    mem[231] = 'd0;
    mem[232] = 'd1020;
    mem[233] = 'd0;
    mem[234] = 'd0;
    mem[235] = 'd1020;
    mem[236] = 'd0;
    mem[237] = 'd1020;
    mem[238] = 'd0;
    mem[239] = 'd0;
    mem[240] = 'd0;
    mem[241] = 'd1020;
    mem[242] = 'd0;
    mem[243] = 'd1020;
    mem[244] = 'd0;
    mem[245] = 'd0;
    mem[246] = 'd0;
    mem[247] = 'd1020;
    mem[248] = 'd0;
    mem[249] = 'd1020;
    mem[250] = 'd0;
    mem[251] = 'd0;
    mem[252] = 'd0;
    mem[253] = 'd1020;
    mem[254] = 'd0;
    mem[255] = 'd1020;
    mem[256] = 'd0;
    mem[257] = 'd0;
    mem[258] = 'd0;
    mem[259] = 'd1020;
    mem[260] = 'd0;
    mem[261] = 'd1020;
    mem[262] = 'd0;
    mem[263] = 'd0;
    mem[264] = 'd0;
    mem[265] = 'd1020;
    mem[266] = 'd0;
    mem[267] = 'd1020;
    mem[268] = 'd0;
    mem[269] = 'd0;
    mem[270] = 'd0;
    mem[271] = 'd1020;
    mem[272] = 'd0;
    mem[273] = 'd1020;
    mem[274] = 'd0;
    mem[275] = 'd0;
    mem[276] = 'd0;
    mem[277] = 'd1020;
    mem[278] = 'd0;
    mem[279] = 'd1020;
    mem[280] = 'd0;
    mem[281] = 'd0;
    mem[282] = 'd0;
    mem[283] = 'd1020;
    mem[284] = 'd0;
    mem[285] = 'd1020;
    mem[286] = 'd0;
    mem[287] = 'd0;
    mem[288] = 'd0;
    mem[289] = 'd1020;
    mem[290] = 'd0;
    mem[291] = 'd1020;
    mem[292] = 'd0;
    mem[293] = 'd0;
    mem[294] = 'd0;
    mem[295] = 'd1020;
    mem[296] = 'd0;
    mem[297] = 'd1020;
    mem[298] = 'd0;
    mem[299] = 'd0;
    mem[300] = 'd0;
    mem[301] = 'd1020;
    mem[302] = 'd0;
    mem[303] = 'd1020;
    mem[304] = 'd0;
    mem[305] = 'd0;
    mem[306] = 'd0;
    mem[307] = 'd1020;
    mem[308] = 'd0;
    mem[309] = 'd1020;
    mem[310] = 'd0;
    mem[311] = 'd0;
    mem[312] = 'd0;
    mem[313] = 'd1020;
    mem[314] = 'd0;
    mem[315] = 'd1020;
    mem[316] = 'd0;
    mem[317] = 'd0;
    mem[318] = 'd0;
    mem[319] = 'd1020;
    mem[320] = 'd0;
    mem[321] = 'd1020;
    mem[322] = 'd0;
    mem[323] = 'd0;
    mem[324] = 'd0;
    mem[325] = 'd1020;
    mem[326] = 'd0;
    mem[327] = 'd1020;
    mem[328] = 'd0;
    mem[329] = 'd0;
    mem[330] = 'd0;
    mem[331] = 'd1020;
    mem[332] = 'd0;
    mem[333] = 'd1020;
    mem[334] = 'd0;
    mem[335] = 'd0;
    mem[336] = 'd0;
    mem[337] = 'd1020;
    mem[338] = 'd0;
    mem[339] = 'd1020;
    mem[340] = 'd0;
    mem[341] = 'd0;
    mem[342] = 'd0;
    mem[343] = 'd1020;
    mem[344] = 'd0;
    mem[345] = 'd1020;
    mem[346] = 'd0;
    mem[347] = 'd0;
    mem[348] = 'd0;
    mem[349] = 'd1020;
    mem[350] = 'd0;
    mem[351] = 'd1020;
    mem[352] = 'd0;
    mem[353] = 'd0;
    mem[354] = 'd0;
    mem[355] = 'd1020;
    mem[356] = 'd0;
    mem[357] = 'd1020;
    mem[358] = 'd0;
    mem[359] = 'd0;
    mem[360] = 'd0;
    mem[361] = 'd1020;
    mem[362] = 'd0;
    mem[363] = 'd1020;
    mem[364] = 'd0;
    mem[365] = 'd0;
    mem[366] = 'd0;
    mem[367] = 'd1020;
    mem[368] = 'd0;
    mem[369] = 'd1020;
    mem[370] = 'd0;
    mem[371] = 'd0;
    mem[372] = 'd0;
    mem[373] = 'd1020;
    mem[374] = 'd0;
    mem[375] = 'd1020;
    mem[376] = 'd0;
    mem[377] = 'd0;
    mem[378] = 'd0;
    mem[379] = 'd1020;
    mem[380] = 'd0;
    mem[381] = 'd1020;
    mem[382] = 'd0;
    mem[383] = 'd0;
    mem[384] = 'd0;
    mem[385] = 'd1020;
    mem[386] = 'd0;
    mem[387] = 'd1020;
    mem[388] = 'd0;
    mem[389] = 'd0;
    mem[390] = 'd0;
    mem[391] = 'd1020;
    mem[392] = 'd0;
    mem[393] = 'd1020;
    mem[394] = 'd0;
    mem[395] = 'd0;
    mem[396] = 'd0;
    mem[397] = 'd1020;
    mem[398] = 'd0;
    mem[399] = 'd1020;
    mem[400] = 'd0;
    mem[401] = 'd0;
    mem[402] = 'd0;
    mem[403] = 'd1020;
    mem[404] = 'd0;
    mem[405] = 'd1020;
    mem[406] = 'd0;
    mem[407] = 'd0;
    mem[408] = 'd0;
    mem[409] = 'd1020;
    mem[410] = 'd0;
    mem[411] = 'd1020;
    mem[412] = 'd0;
    mem[413] = 'd0;
    mem[414] = 'd0;
    mem[415] = 'd1020;
    mem[416] = 'd0;
    mem[417] = 'd1020;
    mem[418] = 'd0;
    mem[419] = 'd0;
    mem[420] = 'd0;
    mem[421] = 'd1020;
    mem[422] = 'd0;
    mem[423] = 'd1020;
    mem[424] = 'd0;
    mem[425] = 'd0;
    mem[426] = 'd0;
    mem[427] = 'd1020;
    mem[428] = 'd0;
    mem[429] = 'd1020;
    mem[430] = 'd0;
    mem[431] = 'd0;
    mem[432] = 'd0;
    mem[433] = 'd1020;
    mem[434] = 'd0;
    mem[435] = 'd1020;
    mem[436] = 'd0;
    mem[437] = 'd0;
    mem[438] = 'd0;
    mem[439] = 'd1020;
    mem[440] = 'd0;
    mem[441] = 'd1020;
    mem[442] = 'd0;
    mem[443] = 'd0;
    mem[444] = 'd0;
    mem[445] = 'd1020;
    mem[446] = 'd0;
    mem[447] = 'd1020;
    mem[448] = 'd0;
    mem[449] = 'd0;
    mem[450] = 'd0;
    mem[451] = 'd1020;
    mem[452] = 'd0;
    mem[453] = 'd1020;
    mem[454] = 'd0;
    mem[455] = 'd0;
    mem[456] = 'd0;
    mem[457] = 'd1020;
    mem[458] = 'd0;
    mem[459] = 'd1020;
    mem[460] = 'd0;
    mem[461] = 'd0;
    mem[462] = 'd0;
    mem[463] = 'd1020;
    mem[464] = 'd0;
    mem[465] = 'd1020;
    mem[466] = 'd0;
    mem[467] = 'd0;
    mem[468] = 'd0;
    mem[469] = 'd0;
    mem[470] = 'd1020;
    mem[471] = 'd0;
    mem[472] = 'd1020;
    mem[473] = 'd0;
    mem[474] = 'd0;
    mem[475] = 'd0;
    mem[476] = 'd1020;
    mem[477] = 'd0;
    mem[478] = 'd1020;
    mem[479] = 'd0;
    mem[480] = 'd0;
    mem[481] = 'd0;
    mem[482] = 'd1020;
    mem[483] = 'd0;
    mem[484] = 'd1020;
    mem[485] = 'd0;
    mem[486] = 'd0;
    mem[487] = 'd0;
    mem[488] = 'd1020;
    mem[489] = 'd0;
    mem[490] = 'd1020;
    mem[491] = 'd0;
    mem[492] = 'd0;
    mem[493] = 'd0;
    mem[494] = 'd1020;
    mem[495] = 'd0;
    mem[496] = 'd1020;
    mem[497] = 'd0;
    mem[498] = 'd0;
    mem[499] = 'd0;
    mem[500] = 'd1020;
    mem[501] = 'd0;
    mem[502] = 'd1020;
    mem[503] = 'd0;
    mem[504] = 'd0;
    mem[505] = 'd0;
    mem[506] = 'd1020;
    mem[507] = 'd0;
    mem[508] = 'd1020;
    mem[509] = 'd0;
    mem[510] = 'd0;
    mem[511] = 'd0;
    mem[512] = 'd1020;
    mem[513] = 'd0;
    mem[514] = 'd1020;
    mem[515] = 'd0;
    mem[516] = 'd0;
    mem[517] = 'd0;
    mem[518] = 'd1020;
    mem[519] = 'd0;
    mem[520] = 'd1020;
    mem[521] = 'd0;
    mem[522] = 'd0;
    mem[523] = 'd0;
    mem[524] = 'd1020;
    mem[525] = 'd0;
    mem[526] = 'd1020;
    mem[527] = 'd0;
    mem[528] = 'd0;
    mem[529] = 'd0;
    mem[530] = 'd1020;
    mem[531] = 'd0;
    mem[532] = 'd1020;
    mem[533] = 'd0;
    mem[534] = 'd0;
    mem[535] = 'd0;
    mem[536] = 'd1020;
    mem[537] = 'd0;
    mem[538] = 'd1020;
    mem[539] = 'd0;
    mem[540] = 'd0;
    mem[541] = 'd0;
    mem[542] = 'd1020;
    mem[543] = 'd0;
    mem[544] = 'd1020;
    mem[545] = 'd0;
    mem[546] = 'd0;
    mem[547] = 'd0;
    mem[548] = 'd988;
    mem[549] = 'd0;
    mem[550] = 'd1000;
    mem[551] = 'd0;
    mem[552] = 'd0;
    mem[553] = 'd0;
    mem[554] = 'd704;
    mem[555] = 'd0;
    mem[556] = 'd872;
    mem[557] = 'd0;
    mem[558] = 'd0;
    mem[559] = 'd0;
    mem[560] = 'd492;
    mem[561] = 'd0;
    mem[562] = 'd804;
    mem[563] = 'd0;
    mem[564] = 'd0;
    mem[565] = 'd0;
    mem[566] = 'd340;
    mem[567] = 'd0;
    mem[568] = 'd768;
    mem[569] = 'd0;
    mem[570] = 'd0;
    mem[571] = 'd0;
    mem[572] = 'd240;
    mem[573] = 'd0;
    mem[574] = 'd748;
    mem[575] = 'd0;
    mem[576] = 'd0;
    mem[577] = 'd0;
    mem[578] = 'd196;
    mem[579] = 'd0;
    mem[580] = 'd740;
    mem[581] = 'd0;
    mem[582] = 'd0;
    mem[583] = 'd0;
    mem[584] = 'd196;
    mem[585] = 'd0;
    mem[586] = 'd740;
    mem[587] = 'd0;
    mem[588] = 'd0;
    mem[589] = 'd0;
    mem[590] = 'd236;
    mem[591] = 'd0;
    mem[592] = 'd744;
    mem[593] = 'd0;
    mem[594] = 'd0;
    mem[595] = 'd0;
    mem[596] = 'd336;
    mem[597] = 'd0;
    mem[598] = 'd764;
    mem[599] = 'd0;
    mem[600] = 'd0;
    mem[601] = 'd0;
    mem[602] = 'd480;
    mem[603] = 'd0;
    mem[604] = 'd800;
    mem[605] = 'd0;
    mem[606] = 'd0;
    mem[607] = 'd0;
    mem[608] = 'd692;
    mem[609] = 'd0;
    mem[610] = 'd868;
    mem[611] = 'd0;
    mem[612] = 'd0;
    mem[613] = 'd0;
    mem[614] = 'd940;
    mem[615] = 'd0;
    mem[616] = 'd976;
    mem[617] = 'd0;
    mem[618] = 'd0;
    mem[619] = 'd0;
    mem[620] = 'd1020;
    mem[621] = 'd0;
    mem[622] = 'd1020;
    mem[623] = 'd0;
    mem[624] = 'd0;
    mem[625] = 'd0;
    mem[626] = 'd1020;
    mem[627] = 'd0;
    mem[628] = 'd1020;
    mem[629] = 'd0;
    mem[630] = 'd0;
    mem[631] = 'd0;
    mem[632] = 'd1020;
    mem[633] = 'd0;
    mem[634] = 'd1020;
    mem[635] = 'd0;
    mem[636] = 'd0;
    mem[637] = 'd0;
    mem[638] = 'd1020;
    mem[639] = 'd0;
    mem[640] = 'd1020;
    mem[641] = 'd0;
    mem[642] = 'd0;
    mem[643] = 'd0;
    mem[644] = 'd1020;
    mem[645] = 'd0;
    mem[646] = 'd1020;
    mem[647] = 'd0;
    mem[648] = 'd0;
    mem[649] = 'd0;
    mem[650] = 'd1020;
    mem[651] = 'd0;
    mem[652] = 'd1020;
    mem[653] = 'd0;
    mem[654] = 'd0;
    mem[655] = 'd0;
    mem[656] = 'd1020;
    mem[657] = 'd0;
    mem[658] = 'd1020;
    mem[659] = 'd0;
    mem[660] = 'd0;
    mem[661] = 'd0;
    mem[662] = 'd1020;
    mem[663] = 'd0;
    mem[664] = 'd1020;
    mem[665] = 'd0;
    mem[666] = 'd0;
    mem[667] = 'd0;
    mem[668] = 'd1020;
    mem[669] = 'd0;
    mem[670] = 'd1020;
    mem[671] = 'd0;
    mem[672] = 'd0;
    mem[673] = 'd0;
    mem[674] = 'd1020;
    mem[675] = 'd0;
    mem[676] = 'd1020;
    mem[677] = 'd0;
    mem[678] = 'd0;
    mem[679] = 'd0;
    mem[680] = 'd1020;
    mem[681] = 'd0;
    mem[682] = 'd1020;
    mem[683] = 'd0;
    mem[684] = 'd0;
    mem[685] = 'd0;
    mem[686] = 'd1020;
    mem[687] = 'd0;
    mem[688] = 'd1020;
    mem[689] = 'd0;
    mem[690] = 'd0;
    mem[691] = 'd0;
    mem[692] = 'd1020;
    mem[693] = 'd0;
    mem[694] = 'd1020;
    mem[695] = 'd0;
    mem[696] = 'd0;
    mem[697] = 'd0;
    mem[698] = 'd1020;
    mem[699] = 'd0;
    mem[700] = 'd1020;
    mem[701] = 'd0;
    mem[702] = 'd0;
    mem[703] = 'd1020;
    mem[704] = 'd0;
    mem[705] = 'd1020;
    mem[706] = 'd0;
    mem[707] = 'd0;
    mem[708] = 'd0;
    mem[709] = 'd1020;
    mem[710] = 'd0;
    mem[711] = 'd1020;
    mem[712] = 'd0;
    mem[713] = 'd0;
    mem[714] = 'd0;
    mem[715] = 'd1020;
    mem[716] = 'd0;
    mem[717] = 'd1020;
    mem[718] = 'd0;
    mem[719] = 'd0;
    mem[720] = 'd0;
    mem[721] = 'd1020;
    mem[722] = 'd0;
    mem[723] = 'd1020;
    mem[724] = 'd0;
    mem[725] = 'd0;
    mem[726] = 'd0;
    mem[727] = 'd1020;
    mem[728] = 'd0;
    mem[729] = 'd1020;
    mem[730] = 'd0;
    mem[731] = 'd0;
    mem[732] = 'd0;
    mem[733] = 'd1020;
    mem[734] = 'd0;
    mem[735] = 'd1020;
    mem[736] = 'd0;
    mem[737] = 'd0;
    mem[738] = 'd0;
    mem[739] = 'd1020;
    mem[740] = 'd0;
    mem[741] = 'd1020;
    mem[742] = 'd0;
    mem[743] = 'd0;
    mem[744] = 'd0;
    mem[745] = 'd1020;
    mem[746] = 'd0;
    mem[747] = 'd1020;
    mem[748] = 'd0;
    mem[749] = 'd0;
    mem[750] = 'd0;
    mem[751] = 'd1020;
    mem[752] = 'd0;
    mem[753] = 'd1020;
    mem[754] = 'd0;
    mem[755] = 'd0;
    mem[756] = 'd0;
    mem[757] = 'd1020;
    mem[758] = 'd0;
    mem[759] = 'd1020;
    mem[760] = 'd0;
    mem[761] = 'd0;
    mem[762] = 'd0;
    mem[763] = 'd1020;
    mem[764] = 'd0;
    mem[765] = 'd1020;
    mem[766] = 'd0;
    mem[767] = 'd0;
    mem[768] = 'd0;
    mem[769] = 'd1020;
    mem[770] = 'd0;
    mem[771] = 'd1020;
    mem[772] = 'd0;
    mem[773] = 'd0;
    mem[774] = 'd0;
    mem[775] = 'd1020;
    mem[776] = 'd0;
    mem[777] = 'd1020;
    mem[778] = 'd0;
    mem[779] = 'd0;
    mem[780] = 'd0;
    mem[781] = 'd1000;
    mem[782] = 'd0;
    mem[783] = 'd1012;
    mem[784] = 'd0;
    mem[785] = 'd0;
    mem[786] = 'd0;
    mem[787] = 'd872;
    mem[788] = 'd0;
    mem[789] = 'd1000;
    mem[790] = 'd0;
    mem[791] = 'd0;
    mem[792] = 'd0;
    mem[793] = 'd804;
    mem[794] = 'd0;
    mem[795] = 'd1000;
    mem[796] = 'd0;
    mem[797] = 'd0;
    mem[798] = 'd0;
    mem[799] = 'd768;
    mem[800] = 'd0;
    mem[801] = 'd1000;
    mem[802] = 'd0;
    mem[803] = 'd0;
    mem[804] = 'd0;
    mem[805] = 'd748;
    mem[806] = 'd0;
    mem[807] = 'd1000;
    mem[808] = 'd0;
    mem[809] = 'd0;
    mem[810] = 'd0;
    mem[811] = 'd740;
    mem[812] = 'd0;
    mem[813] = 'd1000;
    mem[814] = 'd0;
    mem[815] = 'd0;
    mem[816] = 'd0;
    mem[817] = 'd740;
    mem[818] = 'd0;
    mem[819] = 'd1000;
    mem[820] = 'd0;
    mem[821] = 'd0;
    mem[822] = 'd0;
    mem[823] = 'd744;
    mem[824] = 'd0;
    mem[825] = 'd1000;
    mem[826] = 'd0;
    mem[827] = 'd0;
    mem[828] = 'd0;
    mem[829] = 'd764;
    mem[830] = 'd0;
    mem[831] = 'd1000;
    mem[832] = 'd0;
    mem[833] = 'd0;
    mem[834] = 'd0;
    mem[835] = 'd800;
    mem[836] = 'd0;
    mem[837] = 'd1000;
    mem[838] = 'd0;
    mem[839] = 'd0;
    mem[840] = 'd0;
    mem[841] = 'd868;
    mem[842] = 'd0;
    mem[843] = 'd996;
    mem[844] = 'd0;
    mem[845] = 'd0;
    mem[846] = 'd0;
    mem[847] = 'd976;
    mem[848] = 'd0;
    mem[849] = 'd1004;
    mem[850] = 'd0;
    mem[851] = 'd0;
    mem[852] = 'd0;
    mem[853] = 'd1020;
    mem[854] = 'd0;
    mem[855] = 'd1020;
    mem[856] = 'd0;
    mem[857] = 'd0;
    mem[858] = 'd0;
    mem[859] = 'd1020;
    mem[860] = 'd0;
    mem[861] = 'd1020;
    mem[862] = 'd0;
    mem[863] = 'd0;
    mem[864] = 'd0;
    mem[865] = 'd1020;
    mem[866] = 'd0;
    mem[867] = 'd1020;
    mem[868] = 'd0;
    mem[869] = 'd0;
    mem[870] = 'd0;
    mem[871] = 'd1020;
    mem[872] = 'd0;
    mem[873] = 'd1020;
    mem[874] = 'd0;
    mem[875] = 'd0;
    mem[876] = 'd0;
    mem[877] = 'd1020;
    mem[878] = 'd0;
    mem[879] = 'd1020;
    mem[880] = 'd0;
    mem[881] = 'd0;
    mem[882] = 'd0;
    mem[883] = 'd1020;
    mem[884] = 'd0;
    mem[885] = 'd1020;
    mem[886] = 'd0;
    mem[887] = 'd0;
    mem[888] = 'd0;
    mem[889] = 'd1020;
    mem[890] = 'd0;
    mem[891] = 'd1020;
    mem[892] = 'd0;
    mem[893] = 'd0;
    mem[894] = 'd0;
    mem[895] = 'd1020;
    mem[896] = 'd0;
    mem[897] = 'd1020;
    mem[898] = 'd0;
    mem[899] = 'd0;
    mem[900] = 'd0;
    mem[901] = 'd1020;
    mem[902] = 'd0;
    mem[903] = 'd1020;
    mem[904] = 'd0;
    mem[905] = 'd0;
    mem[906] = 'd0;
    mem[907] = 'd1020;
    mem[908] = 'd0;
    mem[909] = 'd1020;
    mem[910] = 'd0;
    mem[911] = 'd0;
    mem[912] = 'd0;
    mem[913] = 'd1020;
    mem[914] = 'd0;
    mem[915] = 'd1020;
    mem[916] = 'd0;
    mem[917] = 'd0;
    mem[918] = 'd0;
    mem[919] = 'd1020;
    mem[920] = 'd0;
    mem[921] = 'd1020;
    mem[922] = 'd0;
    mem[923] = 'd0;
    mem[924] = 'd0;
    mem[925] = 'd1020;
    mem[926] = 'd0;
    mem[927] = 'd1020;
    mem[928] = 'd0;
    mem[929] = 'd0;
    mem[930] = 'd0;
    mem[931] = 'd1020;
    mem[932] = 'd0;
    mem[933] = 'd1020;
    mem[934] = 'd0;
    mem[935] = 'd0;
    mem[936] = 'd0;
    mem[937] = 'd0;
    mem[938] = 'd1020;
    mem[939] = 'd0;
    mem[940] = 'd1020;
    mem[941] = 'd0;
    mem[942] = 'd0;
    mem[943] = 'd0;
    mem[944] = 'd1020;
    mem[945] = 'd0;
    mem[946] = 'd1020;
    mem[947] = 'd0;
    mem[948] = 'd0;
    mem[949] = 'd0;
    mem[950] = 'd1020;
    mem[951] = 'd0;
    mem[952] = 'd1020;
    mem[953] = 'd0;
    mem[954] = 'd0;
    mem[955] = 'd0;
    mem[956] = 'd1020;
    mem[957] = 'd0;
    mem[958] = 'd1020;
    mem[959] = 'd0;
    mem[960] = 'd0;
    mem[961] = 'd0;
    mem[962] = 'd1020;
    mem[963] = 'd0;
    mem[964] = 'd1020;
    mem[965] = 'd0;
    mem[966] = 'd0;
    mem[967] = 'd0;
    mem[968] = 'd1020;
    mem[969] = 'd0;
    mem[970] = 'd1020;
    mem[971] = 'd0;
    mem[972] = 'd0;
    mem[973] = 'd0;
    mem[974] = 'd1020;
    mem[975] = 'd0;
    mem[976] = 'd1020;
    mem[977] = 'd0;
    mem[978] = 'd0;
    mem[979] = 'd0;
    mem[980] = 'd1020;
    mem[981] = 'd0;
    mem[982] = 'd1020;
    mem[983] = 'd0;
    mem[984] = 'd0;
    mem[985] = 'd0;
    mem[986] = 'd1020;
    mem[987] = 'd0;
    mem[988] = 'd1020;
    mem[989] = 'd0;
    mem[990] = 'd0;
    mem[991] = 'd0;
    mem[992] = 'd1020;
    mem[993] = 'd0;
    mem[994] = 'd1020;
    mem[995] = 'd0;
    mem[996] = 'd0;
    mem[997] = 'd0;
    mem[998] = 'd1020;
    mem[999] = 'd0;
    mem[1000] = 'd1020;
    mem[1001] = 'd0;
    mem[1002] = 'd0;
    mem[1003] = 'd0;
    mem[1004] = 'd808;
    mem[1005] = 'd0;
    mem[1006] = 'd912;
    mem[1007] = 'd0;
    mem[1008] = 'd0;
    mem[1009] = 'd0;
    mem[1010] = 'd408;
    mem[1011] = 'd0;
    mem[1012] = 'd768;
    mem[1013] = 'd0;
    mem[1014] = 'd0;
    mem[1015] = 'd0;
    mem[1016] = 'd100;
    mem[1017] = 'd0;
    mem[1018] = 'd696;
    mem[1019] = 'd0;
    mem[1020] = 'd0;
    mem[1021] = 'd0;
    mem[1022] = 'd88;
    mem[1023] = 'd0;
    mem[1024] = 'd772;
    mem[1025] = 'd0;
    mem[1026] = 'd0;
    mem[1027] = 'd0;
    mem[1028] = 'd96;
    mem[1029] = 'd0;
    mem[1030] = 'd828;
    mem[1031] = 'd0;
    mem[1032] = 'd0;
    mem[1033] = 'd0;
    mem[1034] = 'd112;
    mem[1035] = 'd0;
    mem[1036] = 'd868;
    mem[1037] = 'd0;
    mem[1038] = 'd0;
    mem[1039] = 'd0;
    mem[1040] = 'd180;
    mem[1041] = 'd0;
    mem[1042] = 'd900;
    mem[1043] = 'd0;
    mem[1044] = 'd0;
    mem[1045] = 'd0;
    mem[1046] = 'd224;
    mem[1047] = 'd0;
    mem[1048] = 'd916;
    mem[1049] = 'd0;
    mem[1050] = 'd0;
    mem[1051] = 'd0;
    mem[1052] = 'd232;
    mem[1053] = 'd0;
    mem[1054] = 'd916;
    mem[1055] = 'd0;
    mem[1056] = 'd0;
    mem[1057] = 'd0;
    mem[1058] = 'd184;
    mem[1059] = 'd0;
    mem[1060] = 'd900;
    mem[1061] = 'd0;
    mem[1062] = 'd0;
    mem[1063] = 'd0;
    mem[1064] = 'd120;
    mem[1065] = 'd0;
    mem[1066] = 'd868;
    mem[1067] = 'd0;
    mem[1068] = 'd0;
    mem[1069] = 'd0;
    mem[1070] = 'd92;
    mem[1071] = 'd0;
    mem[1072] = 'd828;
    mem[1073] = 'd0;
    mem[1074] = 'd0;
    mem[1075] = 'd0;
    mem[1076] = 'd88;
    mem[1077] = 'd0;
    mem[1078] = 'd776;
    mem[1079] = 'd0;
    mem[1080] = 'd0;
    mem[1081] = 'd0;
    mem[1082] = 'd128;
    mem[1083] = 'd0;
    mem[1084] = 'd712;
    mem[1085] = 'd0;
    mem[1086] = 'd0;
    mem[1087] = 'd0;
    mem[1088] = 'd372;
    mem[1089] = 'd0;
    mem[1090] = 'd752;
    mem[1091] = 'd0;
    mem[1092] = 'd0;
    mem[1093] = 'd0;
    mem[1094] = 'd780;
    mem[1095] = 'd0;
    mem[1096] = 'd904;
    mem[1097] = 'd0;
    mem[1098] = 'd0;
    mem[1099] = 'd0;
    mem[1100] = 'd1012;
    mem[1101] = 'd0;
    mem[1102] = 'd1012;
    mem[1103] = 'd0;
    mem[1104] = 'd0;
    mem[1105] = 'd0;
    mem[1106] = 'd1020;
    mem[1107] = 'd0;
    mem[1108] = 'd1020;
    mem[1109] = 'd0;
    mem[1110] = 'd0;
    mem[1111] = 'd0;
    mem[1112] = 'd1020;
    mem[1113] = 'd0;
    mem[1114] = 'd1020;
    mem[1115] = 'd0;
    mem[1116] = 'd0;
    mem[1117] = 'd0;
    mem[1118] = 'd1020;
    mem[1119] = 'd0;
    mem[1120] = 'd1020;
    mem[1121] = 'd0;
    mem[1122] = 'd0;
    mem[1123] = 'd0;
    mem[1124] = 'd1020;
    mem[1125] = 'd0;
    mem[1126] = 'd1020;
    mem[1127] = 'd0;
    mem[1128] = 'd0;
    mem[1129] = 'd0;
    mem[1130] = 'd1020;
    mem[1131] = 'd0;
    mem[1132] = 'd1020;
    mem[1133] = 'd0;
    mem[1134] = 'd0;
    mem[1135] = 'd0;
    mem[1136] = 'd1020;
    mem[1137] = 'd0;
    mem[1138] = 'd1020;
    mem[1139] = 'd0;
    mem[1140] = 'd0;
    mem[1141] = 'd0;
    mem[1142] = 'd1020;
    mem[1143] = 'd0;
    mem[1144] = 'd1020;
    mem[1145] = 'd0;
    mem[1146] = 'd0;
    mem[1147] = 'd0;
    mem[1148] = 'd1020;
    mem[1149] = 'd0;
    mem[1150] = 'd1020;
    mem[1151] = 'd0;
    mem[1152] = 'd0;
    mem[1153] = 'd0;
    mem[1154] = 'd1020;
    mem[1155] = 'd0;
    mem[1156] = 'd1020;
    mem[1157] = 'd0;
    mem[1158] = 'd0;
    mem[1159] = 'd0;
    mem[1160] = 'd1020;
    mem[1161] = 'd0;
    mem[1162] = 'd1020;
    mem[1163] = 'd0;
    mem[1164] = 'd0;
    mem[1165] = 'd0;
    mem[1166] = 'd1020;
    mem[1167] = 'd0;
    mem[1168] = 'd1020;
    mem[1169] = 'd0;
    mem[1170] = 'd0;
    mem[1171] = 'd1020;
    mem[1172] = 'd0;
    mem[1173] = 'd1020;
    mem[1174] = 'd0;
    mem[1175] = 'd0;
    mem[1176] = 'd0;
    mem[1177] = 'd1020;
    mem[1178] = 'd0;
    mem[1179] = 'd1020;
    mem[1180] = 'd0;
    mem[1181] = 'd0;
    mem[1182] = 'd0;
    mem[1183] = 'd1020;
    mem[1184] = 'd0;
    mem[1185] = 'd1020;
    mem[1186] = 'd0;
    mem[1187] = 'd0;
    mem[1188] = 'd0;
    mem[1189] = 'd1020;
    mem[1190] = 'd0;
    mem[1191] = 'd1020;
    mem[1192] = 'd0;
    mem[1193] = 'd0;
    mem[1194] = 'd0;
    mem[1195] = 'd1020;
    mem[1196] = 'd0;
    mem[1197] = 'd1020;
    mem[1198] = 'd0;
    mem[1199] = 'd0;
    mem[1200] = 'd0;
    mem[1201] = 'd1020;
    mem[1202] = 'd0;
    mem[1203] = 'd1020;
    mem[1204] = 'd0;
    mem[1205] = 'd0;
    mem[1206] = 'd0;
    mem[1207] = 'd1020;
    mem[1208] = 'd0;
    mem[1209] = 'd1020;
    mem[1210] = 'd0;
    mem[1211] = 'd0;
    mem[1212] = 'd0;
    mem[1213] = 'd1020;
    mem[1214] = 'd0;
    mem[1215] = 'd1020;
    mem[1216] = 'd0;
    mem[1217] = 'd0;
    mem[1218] = 'd0;
    mem[1219] = 'd1020;
    mem[1220] = 'd0;
    mem[1221] = 'd1020;
    mem[1222] = 'd0;
    mem[1223] = 'd0;
    mem[1224] = 'd0;
    mem[1225] = 'd1020;
    mem[1226] = 'd0;
    mem[1227] = 'd1020;
    mem[1228] = 'd0;
    mem[1229] = 'd0;
    mem[1230] = 'd0;
    mem[1231] = 'd1020;
    mem[1232] = 'd0;
    mem[1233] = 'd1020;
    mem[1234] = 'd0;
    mem[1235] = 'd0;
    mem[1236] = 'd0;
    mem[1237] = 'd912;
    mem[1238] = 'd0;
    mem[1239] = 'd996;
    mem[1240] = 'd0;
    mem[1241] = 'd0;
    mem[1242] = 'd0;
    mem[1243] = 'd768;
    mem[1244] = 'd0;
    mem[1245] = 'd996;
    mem[1246] = 'd0;
    mem[1247] = 'd0;
    mem[1248] = 'd0;
    mem[1249] = 'd696;
    mem[1250] = 'd0;
    mem[1251] = 'd1012;
    mem[1252] = 'd0;
    mem[1253] = 'd0;
    mem[1254] = 'd0;
    mem[1255] = 'd772;
    mem[1256] = 'd0;
    mem[1257] = 'd1020;
    mem[1258] = 'd0;
    mem[1259] = 'd0;
    mem[1260] = 'd0;
    mem[1261] = 'd828;
    mem[1262] = 'd0;
    mem[1263] = 'd1020;
    mem[1264] = 'd0;
    mem[1265] = 'd0;
    mem[1266] = 'd0;
    mem[1267] = 'd868;
    mem[1268] = 'd0;
    mem[1269] = 'd1020;
    mem[1270] = 'd0;
    mem[1271] = 'd0;
    mem[1272] = 'd0;
    mem[1273] = 'd900;
    mem[1274] = 'd0;
    mem[1275] = 'd1020;
    mem[1276] = 'd0;
    mem[1277] = 'd0;
    mem[1278] = 'd0;
    mem[1279] = 'd916;
    mem[1280] = 'd0;
    mem[1281] = 'd1020;
    mem[1282] = 'd0;
    mem[1283] = 'd0;
    mem[1284] = 'd0;
    mem[1285] = 'd916;
    mem[1286] = 'd0;
    mem[1287] = 'd1020;
    mem[1288] = 'd0;
    mem[1289] = 'd0;
    mem[1290] = 'd0;
    mem[1291] = 'd900;
    mem[1292] = 'd0;
    mem[1293] = 'd1020;
    mem[1294] = 'd0;
    mem[1295] = 'd0;
    mem[1296] = 'd0;
    mem[1297] = 'd868;
    mem[1298] = 'd0;
    mem[1299] = 'd1020;
    mem[1300] = 'd0;
    mem[1301] = 'd0;
    mem[1302] = 'd0;
    mem[1303] = 'd828;
    mem[1304] = 'd0;
    mem[1305] = 'd1020;
    mem[1306] = 'd0;
    mem[1307] = 'd0;
    mem[1308] = 'd0;
    mem[1309] = 'd776;
    mem[1310] = 'd0;
    mem[1311] = 'd1020;
    mem[1312] = 'd0;
    mem[1313] = 'd0;
    mem[1314] = 'd0;
    mem[1315] = 'd712;
    mem[1316] = 'd0;
    mem[1317] = 'd1008;
    mem[1318] = 'd0;
    mem[1319] = 'd0;
    mem[1320] = 'd0;
    mem[1321] = 'd752;
    mem[1322] = 'd0;
    mem[1323] = 'd996;
    mem[1324] = 'd0;
    mem[1325] = 'd0;
    mem[1326] = 'd0;
    mem[1327] = 'd904;
    mem[1328] = 'd0;
    mem[1329] = 'd1000;
    mem[1330] = 'd0;
    mem[1331] = 'd0;
    mem[1332] = 'd0;
    mem[1333] = 'd1012;
    mem[1334] = 'd0;
    mem[1335] = 'd1016;
    mem[1336] = 'd0;
    mem[1337] = 'd0;
    mem[1338] = 'd0;
    mem[1339] = 'd1020;
    mem[1340] = 'd0;
    mem[1341] = 'd1020;
    mem[1342] = 'd0;
    mem[1343] = 'd0;
    mem[1344] = 'd0;
    mem[1345] = 'd1020;
    mem[1346] = 'd0;
    mem[1347] = 'd1020;
    mem[1348] = 'd0;
    mem[1349] = 'd0;
    mem[1350] = 'd0;
    mem[1351] = 'd1020;
    mem[1352] = 'd0;
    mem[1353] = 'd1020;
    mem[1354] = 'd0;
    mem[1355] = 'd0;
    mem[1356] = 'd0;
    mem[1357] = 'd1020;
    mem[1358] = 'd0;
    mem[1359] = 'd1020;
    mem[1360] = 'd0;
    mem[1361] = 'd0;
    mem[1362] = 'd0;
    mem[1363] = 'd1020;
    mem[1364] = 'd0;
    mem[1365] = 'd1020;
    mem[1366] = 'd0;
    mem[1367] = 'd0;
    mem[1368] = 'd0;
    mem[1369] = 'd1020;
    mem[1370] = 'd0;
    mem[1371] = 'd1020;
    mem[1372] = 'd0;
    mem[1373] = 'd0;
    mem[1374] = 'd0;
    mem[1375] = 'd1020;
    mem[1376] = 'd0;
    mem[1377] = 'd1020;
    mem[1378] = 'd0;
    mem[1379] = 'd0;
    mem[1380] = 'd0;
    mem[1381] = 'd1020;
    mem[1382] = 'd0;
    mem[1383] = 'd1020;
    mem[1384] = 'd0;
    mem[1385] = 'd0;
    mem[1386] = 'd0;
    mem[1387] = 'd1020;
    mem[1388] = 'd0;
    mem[1389] = 'd1020;
    mem[1390] = 'd0;
    mem[1391] = 'd0;
    mem[1392] = 'd0;
    mem[1393] = 'd1020;
    mem[1394] = 'd0;
    mem[1395] = 'd1020;
    mem[1396] = 'd0;
    mem[1397] = 'd0;
    mem[1398] = 'd0;
    mem[1399] = 'd1020;
    mem[1400] = 'd0;
    mem[1401] = 'd1020;
    mem[1402] = 'd0;
    mem[1403] = 'd0;
    mem[1404] = 'd0;
    mem[1405] = 'd0;
    mem[1406] = 'd1020;
    mem[1407] = 'd0;
    mem[1408] = 'd1020;
    mem[1409] = 'd0;
    mem[1410] = 'd0;
    mem[1411] = 'd0;
    mem[1412] = 'd1020;
    mem[1413] = 'd0;
    mem[1414] = 'd1020;
    mem[1415] = 'd0;
    mem[1416] = 'd0;
    mem[1417] = 'd0;
    mem[1418] = 'd1020;
    mem[1419] = 'd0;
    mem[1420] = 'd1020;
    mem[1421] = 'd0;
    mem[1422] = 'd0;
    mem[1423] = 'd0;
    mem[1424] = 'd1020;
    mem[1425] = 'd0;
    mem[1426] = 'd1020;
    mem[1427] = 'd0;
    mem[1428] = 'd0;
    mem[1429] = 'd0;
    mem[1430] = 'd1020;
    mem[1431] = 'd0;
    mem[1432] = 'd1020;
    mem[1433] = 'd0;
    mem[1434] = 'd0;
    mem[1435] = 'd0;
    mem[1436] = 'd1020;
    mem[1437] = 'd0;
    mem[1438] = 'd1020;
    mem[1439] = 'd0;
    mem[1440] = 'd0;
    mem[1441] = 'd0;
    mem[1442] = 'd1020;
    mem[1443] = 'd0;
    mem[1444] = 'd1020;
    mem[1445] = 'd0;
    mem[1446] = 'd0;
    mem[1447] = 'd0;
    mem[1448] = 'd1020;
    mem[1449] = 'd0;
    mem[1450] = 'd1020;
    mem[1451] = 'd0;
    mem[1452] = 'd0;
    mem[1453] = 'd0;
    mem[1454] = 'd1020;
    mem[1455] = 'd0;
    mem[1456] = 'd1020;
    mem[1457] = 'd0;
    mem[1458] = 'd0;
    mem[1459] = 'd0;
    mem[1460] = 'd868;
    mem[1461] = 'd0;
    mem[1462] = 'd936;
    mem[1463] = 'd0;
    mem[1464] = 'd0;
    mem[1465] = 'd0;
    mem[1466] = 'd316;
    mem[1467] = 'd0;
    mem[1468] = 'd724;
    mem[1469] = 'd0;
    mem[1470] = 'd0;
    mem[1471] = 'd0;
    mem[1472] = 'd52;
    mem[1473] = 'd0;
    mem[1474] = 'd704;
    mem[1475] = 'd0;
    mem[1476] = 'd0;
    mem[1477] = 'd0;
    mem[1478] = 'd68;
    mem[1479] = 'd0;
    mem[1480] = 'd792;
    mem[1481] = 'd0;
    mem[1482] = 'd0;
    mem[1483] = 'd0;
    mem[1484] = 'd164;
    mem[1485] = 'd0;
    mem[1486] = 'd872;
    mem[1487] = 'd0;
    mem[1488] = 'd0;
    mem[1489] = 'd0;
    mem[1490] = 'd480;
    mem[1491] = 'd0;
    mem[1492] = 'd952;
    mem[1493] = 'd0;
    mem[1494] = 'd0;
    mem[1495] = 'd0;
    mem[1496] = 'd704;
    mem[1497] = 'd0;
    mem[1498] = 'd992;
    mem[1499] = 'd0;
    mem[1500] = 'd0;
    mem[1501] = 'd0;
    mem[1502] = 'd868;
    mem[1503] = 'd0;
    mem[1504] = 'd1012;
    mem[1505] = 'd0;
    mem[1506] = 'd0;
    mem[1507] = 'd0;
    mem[1508] = 'd924;
    mem[1509] = 'd0;
    mem[1510] = 'd1016;
    mem[1511] = 'd0;
    mem[1512] = 'd0;
    mem[1513] = 'd0;
    mem[1514] = 'd940;
    mem[1515] = 'd0;
    mem[1516] = 'd1016;
    mem[1517] = 'd0;
    mem[1518] = 'd0;
    mem[1519] = 'd0;
    mem[1520] = 'd940;
    mem[1521] = 'd0;
    mem[1522] = 'd1016;
    mem[1523] = 'd0;
    mem[1524] = 'd0;
    mem[1525] = 'd0;
    mem[1526] = 'd928;
    mem[1527] = 'd0;
    mem[1528] = 'd1016;
    mem[1529] = 'd0;
    mem[1530] = 'd0;
    mem[1531] = 'd0;
    mem[1532] = 'd876;
    mem[1533] = 'd0;
    mem[1534] = 'd1012;
    mem[1535] = 'd0;
    mem[1536] = 'd0;
    mem[1537] = 'd0;
    mem[1538] = 'd736;
    mem[1539] = 'd0;
    mem[1540] = 'd992;
    mem[1541] = 'd0;
    mem[1542] = 'd0;
    mem[1543] = 'd0;
    mem[1544] = 'd516;
    mem[1545] = 'd0;
    mem[1546] = 'd956;
    mem[1547] = 'd0;
    mem[1548] = 'd0;
    mem[1549] = 'd0;
    mem[1550] = 'd228;
    mem[1551] = 'd0;
    mem[1552] = 'd876;
    mem[1553] = 'd0;
    mem[1554] = 'd0;
    mem[1555] = 'd0;
    mem[1556] = 'd72;
    mem[1557] = 'd0;
    mem[1558] = 'd792;
    mem[1559] = 'd0;
    mem[1560] = 'd0;
    mem[1561] = 'd0;
    mem[1562] = 'd64;
    mem[1563] = 'd0;
    mem[1564] = 'd708;
    mem[1565] = 'd0;
    mem[1566] = 'd0;
    mem[1567] = 'd0;
    mem[1568] = 'd308;
    mem[1569] = 'd0;
    mem[1570] = 'd724;
    mem[1571] = 'd0;
    mem[1572] = 'd0;
    mem[1573] = 'd0;
    mem[1574] = 'd824;
    mem[1575] = 'd0;
    mem[1576] = 'd924;
    mem[1577] = 'd0;
    mem[1578] = 'd0;
    mem[1579] = 'd0;
    mem[1580] = 'd1020;
    mem[1581] = 'd0;
    mem[1582] = 'd1020;
    mem[1583] = 'd0;
    mem[1584] = 'd0;
    mem[1585] = 'd0;
    mem[1586] = 'd1020;
    mem[1587] = 'd0;
    mem[1588] = 'd1020;
    mem[1589] = 'd0;
    mem[1590] = 'd0;
    mem[1591] = 'd0;
    mem[1592] = 'd1020;
    mem[1593] = 'd0;
    mem[1594] = 'd1020;
    mem[1595] = 'd0;
    mem[1596] = 'd0;
    mem[1597] = 'd0;
    mem[1598] = 'd1020;
    mem[1599] = 'd0;
    mem[1600] = 'd1020;
    mem[1601] = 'd0;
    mem[1602] = 'd0;
    mem[1603] = 'd0;
    mem[1604] = 'd1020;
    mem[1605] = 'd0;
    mem[1606] = 'd1020;
    mem[1607] = 'd0;
    mem[1608] = 'd0;
    mem[1609] = 'd0;
    mem[1610] = 'd1020;
    mem[1611] = 'd0;
    mem[1612] = 'd1020;
    mem[1613] = 'd0;
    mem[1614] = 'd0;
    mem[1615] = 'd0;
    mem[1616] = 'd1020;
    mem[1617] = 'd0;
    mem[1618] = 'd1020;
    mem[1619] = 'd0;
    mem[1620] = 'd0;
    mem[1621] = 'd0;
    mem[1622] = 'd1020;
    mem[1623] = 'd0;
    mem[1624] = 'd1020;
    mem[1625] = 'd0;
    mem[1626] = 'd0;
    mem[1627] = 'd0;
    mem[1628] = 'd1020;
    mem[1629] = 'd0;
    mem[1630] = 'd1020;
    mem[1631] = 'd0;
    mem[1632] = 'd0;
    mem[1633] = 'd0;
    mem[1634] = 'd1020;
    mem[1635] = 'd0;
    mem[1636] = 'd1020;
    mem[1637] = 'd0;
    mem[1638] = 'd0;
    mem[1639] = 'd1020;
    mem[1640] = 'd0;
    mem[1641] = 'd1020;
    mem[1642] = 'd0;
    mem[1643] = 'd0;
    mem[1644] = 'd0;
    mem[1645] = 'd1020;
    mem[1646] = 'd0;
    mem[1647] = 'd1020;
    mem[1648] = 'd0;
    mem[1649] = 'd0;
    mem[1650] = 'd0;
    mem[1651] = 'd1020;
    mem[1652] = 'd0;
    mem[1653] = 'd1020;
    mem[1654] = 'd0;
    mem[1655] = 'd0;
    mem[1656] = 'd0;
    mem[1657] = 'd1020;
    mem[1658] = 'd0;
    mem[1659] = 'd1020;
    mem[1660] = 'd0;
    mem[1661] = 'd0;
    mem[1662] = 'd0;
    mem[1663] = 'd1020;
    mem[1664] = 'd0;
    mem[1665] = 'd1020;
    mem[1666] = 'd0;
    mem[1667] = 'd0;
    mem[1668] = 'd0;
    mem[1669] = 'd1020;
    mem[1670] = 'd0;
    mem[1671] = 'd1020;
    mem[1672] = 'd0;
    mem[1673] = 'd0;
    mem[1674] = 'd0;
    mem[1675] = 'd1020;
    mem[1676] = 'd0;
    mem[1677] = 'd1020;
    mem[1678] = 'd0;
    mem[1679] = 'd0;
    mem[1680] = 'd0;
    mem[1681] = 'd1020;
    mem[1682] = 'd0;
    mem[1683] = 'd1020;
    mem[1684] = 'd0;
    mem[1685] = 'd0;
    mem[1686] = 'd0;
    mem[1687] = 'd1020;
    mem[1688] = 'd0;
    mem[1689] = 'd1020;
    mem[1690] = 'd0;
    mem[1691] = 'd0;
    mem[1692] = 'd0;
    mem[1693] = 'd936;
    mem[1694] = 'd0;
    mem[1695] = 'd996;
    mem[1696] = 'd0;
    mem[1697] = 'd0;
    mem[1698] = 'd0;
    mem[1699] = 'd724;
    mem[1700] = 'd0;
    mem[1701] = 'd996;
    mem[1702] = 'd0;
    mem[1703] = 'd0;
    mem[1704] = 'd0;
    mem[1705] = 'd704;
    mem[1706] = 'd0;
    mem[1707] = 'd1020;
    mem[1708] = 'd0;
    mem[1709] = 'd0;
    mem[1710] = 'd0;
    mem[1711] = 'd792;
    mem[1712] = 'd0;
    mem[1713] = 'd1020;
    mem[1714] = 'd0;
    mem[1715] = 'd0;
    mem[1716] = 'd0;
    mem[1717] = 'd872;
    mem[1718] = 'd0;
    mem[1719] = 'd1020;
    mem[1720] = 'd0;
    mem[1721] = 'd0;
    mem[1722] = 'd0;
    mem[1723] = 'd952;
    mem[1724] = 'd0;
    mem[1725] = 'd1020;
    mem[1726] = 'd0;
    mem[1727] = 'd0;
    mem[1728] = 'd0;
    mem[1729] = 'd992;
    mem[1730] = 'd0;
    mem[1731] = 'd1020;
    mem[1732] = 'd0;
    mem[1733] = 'd0;
    mem[1734] = 'd0;
    mem[1735] = 'd1012;
    mem[1736] = 'd0;
    mem[1737] = 'd1020;
    mem[1738] = 'd0;
    mem[1739] = 'd0;
    mem[1740] = 'd0;
    mem[1741] = 'd1016;
    mem[1742] = 'd0;
    mem[1743] = 'd1020;
    mem[1744] = 'd0;
    mem[1745] = 'd0;
    mem[1746] = 'd0;
    mem[1747] = 'd1016;
    mem[1748] = 'd0;
    mem[1749] = 'd1020;
    mem[1750] = 'd0;
    mem[1751] = 'd0;
    mem[1752] = 'd0;
    mem[1753] = 'd1016;
    mem[1754] = 'd0;
    mem[1755] = 'd1020;
    mem[1756] = 'd0;
    mem[1757] = 'd0;
    mem[1758] = 'd0;
    mem[1759] = 'd1016;
    mem[1760] = 'd0;
    mem[1761] = 'd1020;
    mem[1762] = 'd0;
    mem[1763] = 'd0;
    mem[1764] = 'd0;
    mem[1765] = 'd1012;
    mem[1766] = 'd0;
    mem[1767] = 'd1020;
    mem[1768] = 'd0;
    mem[1769] = 'd0;
    mem[1770] = 'd0;
    mem[1771] = 'd992;
    mem[1772] = 'd0;
    mem[1773] = 'd1020;
    mem[1774] = 'd0;
    mem[1775] = 'd0;
    mem[1776] = 'd0;
    mem[1777] = 'd956;
    mem[1778] = 'd0;
    mem[1779] = 'd1020;
    mem[1780] = 'd0;
    mem[1781] = 'd0;
    mem[1782] = 'd0;
    mem[1783] = 'd876;
    mem[1784] = 'd0;
    mem[1785] = 'd1020;
    mem[1786] = 'd0;
    mem[1787] = 'd0;
    mem[1788] = 'd0;
    mem[1789] = 'd792;
    mem[1790] = 'd0;
    mem[1791] = 'd1020;
    mem[1792] = 'd0;
    mem[1793] = 'd0;
    mem[1794] = 'd0;
    mem[1795] = 'd708;
    mem[1796] = 'd0;
    mem[1797] = 'd1016;
    mem[1798] = 'd0;
    mem[1799] = 'd0;
    mem[1800] = 'd0;
    mem[1801] = 'd724;
    mem[1802] = 'd0;
    mem[1803] = 'd996;
    mem[1804] = 'd0;
    mem[1805] = 'd0;
    mem[1806] = 'd0;
    mem[1807] = 'd924;
    mem[1808] = 'd0;
    mem[1809] = 'd1000;
    mem[1810] = 'd0;
    mem[1811] = 'd0;
    mem[1812] = 'd0;
    mem[1813] = 'd1020;
    mem[1814] = 'd0;
    mem[1815] = 'd1020;
    mem[1816] = 'd0;
    mem[1817] = 'd0;
    mem[1818] = 'd0;
    mem[1819] = 'd1020;
    mem[1820] = 'd0;
    mem[1821] = 'd1020;
    mem[1822] = 'd0;
    mem[1823] = 'd0;
    mem[1824] = 'd0;
    mem[1825] = 'd1020;
    mem[1826] = 'd0;
    mem[1827] = 'd1020;
    mem[1828] = 'd0;
    mem[1829] = 'd0;
    mem[1830] = 'd0;
    mem[1831] = 'd1020;
    mem[1832] = 'd0;
    mem[1833] = 'd1020;
    mem[1834] = 'd0;
    mem[1835] = 'd0;
    mem[1836] = 'd0;
    mem[1837] = 'd1020;
    mem[1838] = 'd0;
    mem[1839] = 'd1020;
    mem[1840] = 'd0;
    mem[1841] = 'd0;
    mem[1842] = 'd0;
    mem[1843] = 'd1020;
    mem[1844] = 'd0;
    mem[1845] = 'd1020;
    mem[1846] = 'd0;
    mem[1847] = 'd0;
    mem[1848] = 'd0;
    mem[1849] = 'd1020;
    mem[1850] = 'd0;
    mem[1851] = 'd1020;
    mem[1852] = 'd0;
    mem[1853] = 'd0;
    mem[1854] = 'd0;
    mem[1855] = 'd1020;
    mem[1856] = 'd0;
    mem[1857] = 'd1020;
    mem[1858] = 'd0;
    mem[1859] = 'd0;
    mem[1860] = 'd0;
    mem[1861] = 'd1020;
    mem[1862] = 'd0;
    mem[1863] = 'd1020;
    mem[1864] = 'd0;
    mem[1865] = 'd0;
    mem[1866] = 'd0;
    mem[1867] = 'd1020;
    mem[1868] = 'd0;
    mem[1869] = 'd1020;
    mem[1870] = 'd0;
    mem[1871] = 'd0;
    mem[1872] = 'd0;
    mem[1873] = 'd0;
    mem[1874] = 'd1020;
    mem[1875] = 'd0;
    mem[1876] = 'd1020;
    mem[1877] = 'd0;
    mem[1878] = 'd0;
    mem[1879] = 'd0;
    mem[1880] = 'd1020;
    mem[1881] = 'd0;
    mem[1882] = 'd1020;
    mem[1883] = 'd0;
    mem[1884] = 'd0;
    mem[1885] = 'd0;
    mem[1886] = 'd1020;
    mem[1887] = 'd0;
    mem[1888] = 'd1020;
    mem[1889] = 'd0;
    mem[1890] = 'd0;
    mem[1891] = 'd0;
    mem[1892] = 'd1020;
    mem[1893] = 'd0;
    mem[1894] = 'd1020;
    mem[1895] = 'd0;
    mem[1896] = 'd0;
    mem[1897] = 'd0;
    mem[1898] = 'd1020;
    mem[1899] = 'd0;
    mem[1900] = 'd1020;
    mem[1901] = 'd0;
    mem[1902] = 'd0;
    mem[1903] = 'd0;
    mem[1904] = 'd1020;
    mem[1905] = 'd0;
    mem[1906] = 'd1020;
    mem[1907] = 'd0;
    mem[1908] = 'd0;
    mem[1909] = 'd0;
    mem[1910] = 'd1020;
    mem[1911] = 'd0;
    mem[1912] = 'd1020;
    mem[1913] = 'd0;
    mem[1914] = 'd0;
    mem[1915] = 'd0;
    mem[1916] = 'd1020;
    mem[1917] = 'd0;
    mem[1918] = 'd1020;
    mem[1919] = 'd0;
    mem[1920] = 'd0;
    mem[1921] = 'd0;
    mem[1922] = 'd572;
    mem[1923] = 'd0;
    mem[1924] = 'd804;
    mem[1925] = 'd0;
    mem[1926] = 'd0;
    mem[1927] = 'd0;
    mem[1928] = 'd52;
    mem[1929] = 'd0;
    mem[1930] = 'd660;
    mem[1931] = 'd0;
    mem[1932] = 'd0;
    mem[1933] = 'd0;
    mem[1934] = 'd52;
    mem[1935] = 'd0;
    mem[1936] = 'd764;
    mem[1937] = 'd0;
    mem[1938] = 'd0;
    mem[1939] = 'd0;
    mem[1940] = 'd212;
    mem[1941] = 'd0;
    mem[1942] = 'd868;
    mem[1943] = 'd0;
    mem[1944] = 'd0;
    mem[1945] = 'd0;
    mem[1946] = 'd600;
    mem[1947] = 'd0;
    mem[1948] = 'd972;
    mem[1949] = 'd0;
    mem[1950] = 'd0;
    mem[1951] = 'd0;
    mem[1952] = 'd840;
    mem[1953] = 'd0;
    mem[1954] = 'd1008;
    mem[1955] = 'd0;
    mem[1956] = 'd0;
    mem[1957] = 'd0;
    mem[1958] = 'd852;
    mem[1959] = 'd0;
    mem[1960] = 'd1012;
    mem[1961] = 'd0;
    mem[1962] = 'd0;
    mem[1963] = 'd0;
    mem[1964] = 'd864;
    mem[1965] = 'd0;
    mem[1966] = 'd1012;
    mem[1967] = 'd0;
    mem[1968] = 'd0;
    mem[1969] = 'd0;
    mem[1970] = 'd880;
    mem[1971] = 'd0;
    mem[1972] = 'd1012;
    mem[1973] = 'd0;
    mem[1974] = 'd0;
    mem[1975] = 'd0;
    mem[1976] = 'd888;
    mem[1977] = 'd0;
    mem[1978] = 'd1012;
    mem[1979] = 'd0;
    mem[1980] = 'd0;
    mem[1981] = 'd0;
    mem[1982] = 'd892;
    mem[1983] = 'd0;
    mem[1984] = 'd1012;
    mem[1985] = 'd0;
    mem[1986] = 'd0;
    mem[1987] = 'd0;
    mem[1988] = 'd892;
    mem[1989] = 'd0;
    mem[1990] = 'd1012;
    mem[1991] = 'd0;
    mem[1992] = 'd0;
    mem[1993] = 'd0;
    mem[1994] = 'd888;
    mem[1995] = 'd0;
    mem[1996] = 'd1012;
    mem[1997] = 'd0;
    mem[1998] = 'd0;
    mem[1999] = 'd0;
    mem[2000] = 'd876;
    mem[2001] = 'd0;
    mem[2002] = 'd1012;
    mem[2003] = 'd0;
    mem[2004] = 'd0;
    mem[2005] = 'd0;
    mem[2006] = 'd864;
    mem[2007] = 'd0;
    mem[2008] = 'd1012;
    mem[2009] = 'd0;
    mem[2010] = 'd0;
    mem[2011] = 'd0;
    mem[2012] = 'd848;
    mem[2013] = 'd0;
    mem[2014] = 'd1012;
    mem[2015] = 'd0;
    mem[2016] = 'd0;
    mem[2017] = 'd0;
    mem[2018] = 'd836;
    mem[2019] = 'd0;
    mem[2020] = 'd1012;
    mem[2021] = 'd0;
    mem[2022] = 'd0;
    mem[2023] = 'd0;
    mem[2024] = 'd648;
    mem[2025] = 'd0;
    mem[2026] = 'd976;
    mem[2027] = 'd0;
    mem[2028] = 'd0;
    mem[2029] = 'd0;
    mem[2030] = 'd276;
    mem[2031] = 'd0;
    mem[2032] = 'd880;
    mem[2033] = 'd0;
    mem[2034] = 'd0;
    mem[2035] = 'd0;
    mem[2036] = 'd60;
    mem[2037] = 'd0;
    mem[2038] = 'd768;
    mem[2039] = 'd0;
    mem[2040] = 'd0;
    mem[2041] = 'd0;
    mem[2042] = 'd84;
    mem[2043] = 'd0;
    mem[2044] = 'd680;
    mem[2045] = 'd0;
    mem[2046] = 'd0;
    mem[2047] = 'd0;
    mem[2048] = 'd532;
    mem[2049] = 'd0;
    mem[2050] = 'd792;
    mem[2051] = 'd0;
    mem[2052] = 'd0;
    mem[2053] = 'd0;
    mem[2054] = 'd988;
    mem[2055] = 'd0;
    mem[2056] = 'd1004;
    mem[2057] = 'd0;
    mem[2058] = 'd0;
    mem[2059] = 'd0;
    mem[2060] = 'd1020;
    mem[2061] = 'd0;
    mem[2062] = 'd1020;
    mem[2063] = 'd0;
    mem[2064] = 'd0;
    mem[2065] = 'd0;
    mem[2066] = 'd1020;
    mem[2067] = 'd0;
    mem[2068] = 'd1020;
    mem[2069] = 'd0;
    mem[2070] = 'd0;
    mem[2071] = 'd0;
    mem[2072] = 'd1020;
    mem[2073] = 'd0;
    mem[2074] = 'd1020;
    mem[2075] = 'd0;
    mem[2076] = 'd0;
    mem[2077] = 'd0;
    mem[2078] = 'd1020;
    mem[2079] = 'd0;
    mem[2080] = 'd1020;
    mem[2081] = 'd0;
    mem[2082] = 'd0;
    mem[2083] = 'd0;
    mem[2084] = 'd1020;
    mem[2085] = 'd0;
    mem[2086] = 'd1020;
    mem[2087] = 'd0;
    mem[2088] = 'd0;
    mem[2089] = 'd0;
    mem[2090] = 'd1020;
    mem[2091] = 'd0;
    mem[2092] = 'd1020;
    mem[2093] = 'd0;
    mem[2094] = 'd0;
    mem[2095] = 'd0;
    mem[2096] = 'd1020;
    mem[2097] = 'd0;
    mem[2098] = 'd1020;
    mem[2099] = 'd0;
    mem[2100] = 'd0;
    mem[2101] = 'd0;
    mem[2102] = 'd1020;
    mem[2103] = 'd0;
    mem[2104] = 'd1020;
    mem[2105] = 'd0;
    mem[2106] = 'd0;
    mem[2107] = 'd1020;
    mem[2108] = 'd0;
    mem[2109] = 'd1020;
    mem[2110] = 'd0;
    mem[2111] = 'd0;
    mem[2112] = 'd0;
    mem[2113] = 'd1020;
    mem[2114] = 'd0;
    mem[2115] = 'd1020;
    mem[2116] = 'd0;
    mem[2117] = 'd0;
    mem[2118] = 'd0;
    mem[2119] = 'd1020;
    mem[2120] = 'd0;
    mem[2121] = 'd1020;
    mem[2122] = 'd0;
    mem[2123] = 'd0;
    mem[2124] = 'd0;
    mem[2125] = 'd1020;
    mem[2126] = 'd0;
    mem[2127] = 'd1020;
    mem[2128] = 'd0;
    mem[2129] = 'd0;
    mem[2130] = 'd0;
    mem[2131] = 'd1020;
    mem[2132] = 'd0;
    mem[2133] = 'd1020;
    mem[2134] = 'd0;
    mem[2135] = 'd0;
    mem[2136] = 'd0;
    mem[2137] = 'd1020;
    mem[2138] = 'd0;
    mem[2139] = 'd1020;
    mem[2140] = 'd0;
    mem[2141] = 'd0;
    mem[2142] = 'd0;
    mem[2143] = 'd1020;
    mem[2144] = 'd0;
    mem[2145] = 'd1020;
    mem[2146] = 'd0;
    mem[2147] = 'd0;
    mem[2148] = 'd0;
    mem[2149] = 'd1020;
    mem[2150] = 'd0;
    mem[2151] = 'd1020;
    mem[2152] = 'd0;
    mem[2153] = 'd0;
    mem[2154] = 'd0;
    mem[2155] = 'd804;
    mem[2156] = 'd0;
    mem[2157] = 'd984;
    mem[2158] = 'd0;
    mem[2159] = 'd0;
    mem[2160] = 'd0;
    mem[2161] = 'd660;
    mem[2162] = 'd0;
    mem[2163] = 'd1012;
    mem[2164] = 'd0;
    mem[2165] = 'd0;
    mem[2166] = 'd0;
    mem[2167] = 'd764;
    mem[2168] = 'd0;
    mem[2169] = 'd1020;
    mem[2170] = 'd0;
    mem[2171] = 'd0;
    mem[2172] = 'd0;
    mem[2173] = 'd868;
    mem[2174] = 'd0;
    mem[2175] = 'd1020;
    mem[2176] = 'd0;
    mem[2177] = 'd0;
    mem[2178] = 'd0;
    mem[2179] = 'd972;
    mem[2180] = 'd0;
    mem[2181] = 'd1020;
    mem[2182] = 'd0;
    mem[2183] = 'd0;
    mem[2184] = 'd0;
    mem[2185] = 'd1008;
    mem[2186] = 'd0;
    mem[2187] = 'd1020;
    mem[2188] = 'd0;
    mem[2189] = 'd0;
    mem[2190] = 'd0;
    mem[2191] = 'd1012;
    mem[2192] = 'd0;
    mem[2193] = 'd1020;
    mem[2194] = 'd0;
    mem[2195] = 'd0;
    mem[2196] = 'd0;
    mem[2197] = 'd1012;
    mem[2198] = 'd0;
    mem[2199] = 'd1020;
    mem[2200] = 'd0;
    mem[2201] = 'd0;
    mem[2202] = 'd0;
    mem[2203] = 'd1012;
    mem[2204] = 'd0;
    mem[2205] = 'd1020;
    mem[2206] = 'd0;
    mem[2207] = 'd0;
    mem[2208] = 'd0;
    mem[2209] = 'd1012;
    mem[2210] = 'd0;
    mem[2211] = 'd1020;
    mem[2212] = 'd0;
    mem[2213] = 'd0;
    mem[2214] = 'd0;
    mem[2215] = 'd1012;
    mem[2216] = 'd0;
    mem[2217] = 'd1020;
    mem[2218] = 'd0;
    mem[2219] = 'd0;
    mem[2220] = 'd0;
    mem[2221] = 'd1012;
    mem[2222] = 'd0;
    mem[2223] = 'd1020;
    mem[2224] = 'd0;
    mem[2225] = 'd0;
    mem[2226] = 'd0;
    mem[2227] = 'd1012;
    mem[2228] = 'd0;
    mem[2229] = 'd1020;
    mem[2230] = 'd0;
    mem[2231] = 'd0;
    mem[2232] = 'd0;
    mem[2233] = 'd1012;
    mem[2234] = 'd0;
    mem[2235] = 'd1020;
    mem[2236] = 'd0;
    mem[2237] = 'd0;
    mem[2238] = 'd0;
    mem[2239] = 'd1012;
    mem[2240] = 'd0;
    mem[2241] = 'd1020;
    mem[2242] = 'd0;
    mem[2243] = 'd0;
    mem[2244] = 'd0;
    mem[2245] = 'd1012;
    mem[2246] = 'd0;
    mem[2247] = 'd1020;
    mem[2248] = 'd0;
    mem[2249] = 'd0;
    mem[2250] = 'd0;
    mem[2251] = 'd1012;
    mem[2252] = 'd0;
    mem[2253] = 'd1020;
    mem[2254] = 'd0;
    mem[2255] = 'd0;
    mem[2256] = 'd0;
    mem[2257] = 'd976;
    mem[2258] = 'd0;
    mem[2259] = 'd1020;
    mem[2260] = 'd0;
    mem[2261] = 'd0;
    mem[2262] = 'd0;
    mem[2263] = 'd880;
    mem[2264] = 'd0;
    mem[2265] = 'd1020;
    mem[2266] = 'd0;
    mem[2267] = 'd0;
    mem[2268] = 'd0;
    mem[2269] = 'd768;
    mem[2270] = 'd0;
    mem[2271] = 'd1020;
    mem[2272] = 'd0;
    mem[2273] = 'd0;
    mem[2274] = 'd0;
    mem[2275] = 'd680;
    mem[2276] = 'd0;
    mem[2277] = 'd1012;
    mem[2278] = 'd0;
    mem[2279] = 'd0;
    mem[2280] = 'd0;
    mem[2281] = 'd792;
    mem[2282] = 'd0;
    mem[2283] = 'd996;
    mem[2284] = 'd0;
    mem[2285] = 'd0;
    mem[2286] = 'd0;
    mem[2287] = 'd1004;
    mem[2288] = 'd0;
    mem[2289] = 'd1012;
    mem[2290] = 'd0;
    mem[2291] = 'd0;
    mem[2292] = 'd0;
    mem[2293] = 'd1020;
    mem[2294] = 'd0;
    mem[2295] = 'd1020;
    mem[2296] = 'd0;
    mem[2297] = 'd0;
    mem[2298] = 'd0;
    mem[2299] = 'd1020;
    mem[2300] = 'd0;
    mem[2301] = 'd1020;
    mem[2302] = 'd0;
    mem[2303] = 'd0;
    mem[2304] = 'd0;
    mem[2305] = 'd1020;
    mem[2306] = 'd0;
    mem[2307] = 'd1020;
    mem[2308] = 'd0;
    mem[2309] = 'd0;
    mem[2310] = 'd0;
    mem[2311] = 'd1020;
    mem[2312] = 'd0;
    mem[2313] = 'd1020;
    mem[2314] = 'd0;
    mem[2315] = 'd0;
    mem[2316] = 'd0;
    mem[2317] = 'd1020;
    mem[2318] = 'd0;
    mem[2319] = 'd1020;
    mem[2320] = 'd0;
    mem[2321] = 'd0;
    mem[2322] = 'd0;
    mem[2323] = 'd1020;
    mem[2324] = 'd0;
    mem[2325] = 'd1020;
    mem[2326] = 'd0;
    mem[2327] = 'd0;
    mem[2328] = 'd0;
    mem[2329] = 'd1020;
    mem[2330] = 'd0;
    mem[2331] = 'd1020;
    mem[2332] = 'd0;
    mem[2333] = 'd0;
    mem[2334] = 'd0;
    mem[2335] = 'd1020;
    mem[2336] = 'd0;
    mem[2337] = 'd1020;
    mem[2338] = 'd0;
    mem[2339] = 'd0;
    mem[2340] = 'd0;
    mem[2341] = 'd0;
    mem[2342] = 'd1020;
    mem[2343] = 'd0;
    mem[2344] = 'd1020;
    mem[2345] = 'd0;
    mem[2346] = 'd0;
    mem[2347] = 'd0;
    mem[2348] = 'd1020;
    mem[2349] = 'd0;
    mem[2350] = 'd1020;
    mem[2351] = 'd0;
    mem[2352] = 'd0;
    mem[2353] = 'd0;
    mem[2354] = 'd1020;
    mem[2355] = 'd0;
    mem[2356] = 'd1020;
    mem[2357] = 'd0;
    mem[2358] = 'd0;
    mem[2359] = 'd0;
    mem[2360] = 'd1020;
    mem[2361] = 'd0;
    mem[2362] = 'd1020;
    mem[2363] = 'd0;
    mem[2364] = 'd0;
    mem[2365] = 'd0;
    mem[2366] = 'd1020;
    mem[2367] = 'd0;
    mem[2368] = 'd1020;
    mem[2369] = 'd0;
    mem[2370] = 'd0;
    mem[2371] = 'd0;
    mem[2372] = 'd1020;
    mem[2373] = 'd0;
    mem[2374] = 'd1020;
    mem[2375] = 'd0;
    mem[2376] = 'd0;
    mem[2377] = 'd0;
    mem[2378] = 'd912;
    mem[2379] = 'd0;
    mem[2380] = 'd964;
    mem[2381] = 'd0;
    mem[2382] = 'd0;
    mem[2383] = 'd0;
    mem[2384] = 'd296;
    mem[2385] = 'd0;
    mem[2386] = 'd700;
    mem[2387] = 'd0;
    mem[2388] = 'd0;
    mem[2389] = 'd0;
    mem[2390] = 'd36;
    mem[2391] = 'd0;
    mem[2392] = 'd696;
    mem[2393] = 'd0;
    mem[2394] = 'd0;
    mem[2395] = 'd0;
    mem[2396] = 'd140;
    mem[2397] = 'd0;
    mem[2398] = 'd816;
    mem[2399] = 'd0;
    mem[2400] = 'd0;
    mem[2401] = 'd0;
    mem[2402] = 'd520;
    mem[2403] = 'd0;
    mem[2404] = 'd948;
    mem[2405] = 'd0;
    mem[2406] = 'd0;
    mem[2407] = 'd0;
    mem[2408] = 'd764;
    mem[2409] = 'd0;
    mem[2410] = 'd1004;
    mem[2411] = 'd0;
    mem[2412] = 'd0;
    mem[2413] = 'd0;
    mem[2414] = 'd776;
    mem[2415] = 'd0;
    mem[2416] = 'd1004;
    mem[2417] = 'd0;
    mem[2418] = 'd0;
    mem[2419] = 'd0;
    mem[2420] = 'd788;
    mem[2421] = 'd0;
    mem[2422] = 'd1008;
    mem[2423] = 'd0;
    mem[2424] = 'd0;
    mem[2425] = 'd0;
    mem[2426] = 'd804;
    mem[2427] = 'd0;
    mem[2428] = 'd1008;
    mem[2429] = 'd0;
    mem[2430] = 'd0;
    mem[2431] = 'd0;
    mem[2432] = 'd820;
    mem[2433] = 'd0;
    mem[2434] = 'd1008;
    mem[2435] = 'd0;
    mem[2436] = 'd0;
    mem[2437] = 'd0;
    mem[2438] = 'd836;
    mem[2439] = 'd0;
    mem[2440] = 'd1008;
    mem[2441] = 'd0;
    mem[2442] = 'd0;
    mem[2443] = 'd0;
    mem[2444] = 'd844;
    mem[2445] = 'd0;
    mem[2446] = 'd1012;
    mem[2447] = 'd0;
    mem[2448] = 'd0;
    mem[2449] = 'd0;
    mem[2450] = 'd848;
    mem[2451] = 'd0;
    mem[2452] = 'd1012;
    mem[2453] = 'd0;
    mem[2454] = 'd0;
    mem[2455] = 'd0;
    mem[2456] = 'd848;
    mem[2457] = 'd0;
    mem[2458] = 'd1012;
    mem[2459] = 'd0;
    mem[2460] = 'd0;
    mem[2461] = 'd0;
    mem[2462] = 'd840;
    mem[2463] = 'd0;
    mem[2464] = 'd1012;
    mem[2465] = 'd0;
    mem[2466] = 'd0;
    mem[2467] = 'd0;
    mem[2468] = 'd832;
    mem[2469] = 'd0;
    mem[2470] = 'd1008;
    mem[2471] = 'd0;
    mem[2472] = 'd0;
    mem[2473] = 'd0;
    mem[2474] = 'd816;
    mem[2475] = 'd0;
    mem[2476] = 'd1008;
    mem[2477] = 'd0;
    mem[2478] = 'd0;
    mem[2479] = 'd0;
    mem[2480] = 'd800;
    mem[2481] = 'd0;
    mem[2482] = 'd1008;
    mem[2483] = 'd0;
    mem[2484] = 'd0;
    mem[2485] = 'd0;
    mem[2486] = 'd784;
    mem[2487] = 'd0;
    mem[2488] = 'd1008;
    mem[2489] = 'd0;
    mem[2490] = 'd0;
    mem[2491] = 'd0;
    mem[2492] = 'd772;
    mem[2493] = 'd0;
    mem[2494] = 'd1004;
    mem[2495] = 'd0;
    mem[2496] = 'd0;
    mem[2497] = 'd0;
    mem[2498] = 'd760;
    mem[2499] = 'd0;
    mem[2500] = 'd1008;
    mem[2501] = 'd0;
    mem[2502] = 'd0;
    mem[2503] = 'd0;
    mem[2504] = 'd588;
    mem[2505] = 'd0;
    mem[2506] = 'd964;
    mem[2507] = 'd0;
    mem[2508] = 'd0;
    mem[2509] = 'd0;
    mem[2510] = 'd184;
    mem[2511] = 'd0;
    mem[2512] = 'd828;
    mem[2513] = 'd0;
    mem[2514] = 'd0;
    mem[2515] = 'd0;
    mem[2516] = 'd36;
    mem[2517] = 'd0;
    mem[2518] = 'd700;
    mem[2519] = 'd0;
    mem[2520] = 'd0;
    mem[2521] = 'd0;
    mem[2522] = 'd268;
    mem[2523] = 'd0;
    mem[2524] = 'd688;
    mem[2525] = 'd0;
    mem[2526] = 'd0;
    mem[2527] = 'd0;
    mem[2528] = 'd904;
    mem[2529] = 'd0;
    mem[2530] = 'd960;
    mem[2531] = 'd0;
    mem[2532] = 'd0;
    mem[2533] = 'd0;
    mem[2534] = 'd1020;
    mem[2535] = 'd0;
    mem[2536] = 'd1020;
    mem[2537] = 'd0;
    mem[2538] = 'd0;
    mem[2539] = 'd0;
    mem[2540] = 'd1020;
    mem[2541] = 'd0;
    mem[2542] = 'd1020;
    mem[2543] = 'd0;
    mem[2544] = 'd0;
    mem[2545] = 'd0;
    mem[2546] = 'd1020;
    mem[2547] = 'd0;
    mem[2548] = 'd1020;
    mem[2549] = 'd0;
    mem[2550] = 'd0;
    mem[2551] = 'd0;
    mem[2552] = 'd1020;
    mem[2553] = 'd0;
    mem[2554] = 'd1020;
    mem[2555] = 'd0;
    mem[2556] = 'd0;
    mem[2557] = 'd0;
    mem[2558] = 'd1020;
    mem[2559] = 'd0;
    mem[2560] = 'd1020;
    mem[2561] = 'd0;
    mem[2562] = 'd0;
    mem[2563] = 'd0;
    mem[2564] = 'd1020;
    mem[2565] = 'd0;
    mem[2566] = 'd1020;
    mem[2567] = 'd0;
    mem[2568] = 'd0;
    mem[2569] = 'd0;
    mem[2570] = 'd1020;
    mem[2571] = 'd0;
    mem[2572] = 'd1020;
    mem[2573] = 'd0;
    mem[2574] = 'd0;
    mem[2575] = 'd1020;
    mem[2576] = 'd0;
    mem[2577] = 'd1020;
    mem[2578] = 'd0;
    mem[2579] = 'd0;
    mem[2580] = 'd0;
    mem[2581] = 'd1020;
    mem[2582] = 'd0;
    mem[2583] = 'd1020;
    mem[2584] = 'd0;
    mem[2585] = 'd0;
    mem[2586] = 'd0;
    mem[2587] = 'd1020;
    mem[2588] = 'd0;
    mem[2589] = 'd1020;
    mem[2590] = 'd0;
    mem[2591] = 'd0;
    mem[2592] = 'd0;
    mem[2593] = 'd1020;
    mem[2594] = 'd0;
    mem[2595] = 'd1020;
    mem[2596] = 'd0;
    mem[2597] = 'd0;
    mem[2598] = 'd0;
    mem[2599] = 'd1020;
    mem[2600] = 'd0;
    mem[2601] = 'd1020;
    mem[2602] = 'd0;
    mem[2603] = 'd0;
    mem[2604] = 'd0;
    mem[2605] = 'd1020;
    mem[2606] = 'd0;
    mem[2607] = 'd1020;
    mem[2608] = 'd0;
    mem[2609] = 'd0;
    mem[2610] = 'd0;
    mem[2611] = 'd964;
    mem[2612] = 'd0;
    mem[2613] = 'd1012;
    mem[2614] = 'd0;
    mem[2615] = 'd0;
    mem[2616] = 'd0;
    mem[2617] = 'd700;
    mem[2618] = 'd0;
    mem[2619] = 'd988;
    mem[2620] = 'd0;
    mem[2621] = 'd0;
    mem[2622] = 'd0;
    mem[2623] = 'd696;
    mem[2624] = 'd0;
    mem[2625] = 'd1020;
    mem[2626] = 'd0;
    mem[2627] = 'd0;
    mem[2628] = 'd0;
    mem[2629] = 'd816;
    mem[2630] = 'd0;
    mem[2631] = 'd1020;
    mem[2632] = 'd0;
    mem[2633] = 'd0;
    mem[2634] = 'd0;
    mem[2635] = 'd948;
    mem[2636] = 'd0;
    mem[2637] = 'd1020;
    mem[2638] = 'd0;
    mem[2639] = 'd0;
    mem[2640] = 'd0;
    mem[2641] = 'd1004;
    mem[2642] = 'd0;
    mem[2643] = 'd1020;
    mem[2644] = 'd0;
    mem[2645] = 'd0;
    mem[2646] = 'd0;
    mem[2647] = 'd1004;
    mem[2648] = 'd0;
    mem[2649] = 'd1020;
    mem[2650] = 'd0;
    mem[2651] = 'd0;
    mem[2652] = 'd0;
    mem[2653] = 'd1008;
    mem[2654] = 'd0;
    mem[2655] = 'd1020;
    mem[2656] = 'd0;
    mem[2657] = 'd0;
    mem[2658] = 'd0;
    mem[2659] = 'd1008;
    mem[2660] = 'd0;
    mem[2661] = 'd1020;
    mem[2662] = 'd0;
    mem[2663] = 'd0;
    mem[2664] = 'd0;
    mem[2665] = 'd1008;
    mem[2666] = 'd0;
    mem[2667] = 'd1020;
    mem[2668] = 'd0;
    mem[2669] = 'd0;
    mem[2670] = 'd0;
    mem[2671] = 'd1008;
    mem[2672] = 'd0;
    mem[2673] = 'd1020;
    mem[2674] = 'd0;
    mem[2675] = 'd0;
    mem[2676] = 'd0;
    mem[2677] = 'd1012;
    mem[2678] = 'd0;
    mem[2679] = 'd1020;
    mem[2680] = 'd0;
    mem[2681] = 'd0;
    mem[2682] = 'd0;
    mem[2683] = 'd1012;
    mem[2684] = 'd0;
    mem[2685] = 'd1020;
    mem[2686] = 'd0;
    mem[2687] = 'd0;
    mem[2688] = 'd0;
    mem[2689] = 'd1012;
    mem[2690] = 'd0;
    mem[2691] = 'd1020;
    mem[2692] = 'd0;
    mem[2693] = 'd0;
    mem[2694] = 'd0;
    mem[2695] = 'd1012;
    mem[2696] = 'd0;
    mem[2697] = 'd1020;
    mem[2698] = 'd0;
    mem[2699] = 'd0;
    mem[2700] = 'd0;
    mem[2701] = 'd1008;
    mem[2702] = 'd0;
    mem[2703] = 'd1020;
    mem[2704] = 'd0;
    mem[2705] = 'd0;
    mem[2706] = 'd0;
    mem[2707] = 'd1008;
    mem[2708] = 'd0;
    mem[2709] = 'd1020;
    mem[2710] = 'd0;
    mem[2711] = 'd0;
    mem[2712] = 'd0;
    mem[2713] = 'd1008;
    mem[2714] = 'd0;
    mem[2715] = 'd1020;
    mem[2716] = 'd0;
    mem[2717] = 'd0;
    mem[2718] = 'd0;
    mem[2719] = 'd1008;
    mem[2720] = 'd0;
    mem[2721] = 'd1020;
    mem[2722] = 'd0;
    mem[2723] = 'd0;
    mem[2724] = 'd0;
    mem[2725] = 'd1004;
    mem[2726] = 'd0;
    mem[2727] = 'd1020;
    mem[2728] = 'd0;
    mem[2729] = 'd0;
    mem[2730] = 'd0;
    mem[2731] = 'd1008;
    mem[2732] = 'd0;
    mem[2733] = 'd1020;
    mem[2734] = 'd0;
    mem[2735] = 'd0;
    mem[2736] = 'd0;
    mem[2737] = 'd964;
    mem[2738] = 'd0;
    mem[2739] = 'd1020;
    mem[2740] = 'd0;
    mem[2741] = 'd0;
    mem[2742] = 'd0;
    mem[2743] = 'd828;
    mem[2744] = 'd0;
    mem[2745] = 'd1020;
    mem[2746] = 'd0;
    mem[2747] = 'd0;
    mem[2748] = 'd0;
    mem[2749] = 'd700;
    mem[2750] = 'd0;
    mem[2751] = 'd1020;
    mem[2752] = 'd0;
    mem[2753] = 'd0;
    mem[2754] = 'd0;
    mem[2755] = 'd688;
    mem[2756] = 'd0;
    mem[2757] = 'd988;
    mem[2758] = 'd0;
    mem[2759] = 'd0;
    mem[2760] = 'd0;
    mem[2761] = 'd960;
    mem[2762] = 'd0;
    mem[2763] = 'd1012;
    mem[2764] = 'd0;
    mem[2765] = 'd0;
    mem[2766] = 'd0;
    mem[2767] = 'd1020;
    mem[2768] = 'd0;
    mem[2769] = 'd1020;
    mem[2770] = 'd0;
    mem[2771] = 'd0;
    mem[2772] = 'd0;
    mem[2773] = 'd1020;
    mem[2774] = 'd0;
    mem[2775] = 'd1020;
    mem[2776] = 'd0;
    mem[2777] = 'd0;
    mem[2778] = 'd0;
    mem[2779] = 'd1020;
    mem[2780] = 'd0;
    mem[2781] = 'd1020;
    mem[2782] = 'd0;
    mem[2783] = 'd0;
    mem[2784] = 'd0;
    mem[2785] = 'd1020;
    mem[2786] = 'd0;
    mem[2787] = 'd1020;
    mem[2788] = 'd0;
    mem[2789] = 'd0;
    mem[2790] = 'd0;
    mem[2791] = 'd1020;
    mem[2792] = 'd0;
    mem[2793] = 'd1020;
    mem[2794] = 'd0;
    mem[2795] = 'd0;
    mem[2796] = 'd0;
    mem[2797] = 'd1020;
    mem[2798] = 'd0;
    mem[2799] = 'd1020;
    mem[2800] = 'd0;
    mem[2801] = 'd0;
    mem[2802] = 'd0;
    mem[2803] = 'd1020;
    mem[2804] = 'd0;
    mem[2805] = 'd1020;
    mem[2806] = 'd0;
    mem[2807] = 'd0;
    mem[2808] = 'd0;
    mem[2809] = 'd0;
    mem[2810] = 'd1020;
    mem[2811] = 'd0;
    mem[2812] = 'd1020;
    mem[2813] = 'd0;
    mem[2814] = 'd0;
    mem[2815] = 'd0;
    mem[2816] = 'd1020;
    mem[2817] = 'd0;
    mem[2818] = 'd1020;
    mem[2819] = 'd0;
    mem[2820] = 'd0;
    mem[2821] = 'd0;
    mem[2822] = 'd1020;
    mem[2823] = 'd0;
    mem[2824] = 'd1020;
    mem[2825] = 'd0;
    mem[2826] = 'd0;
    mem[2827] = 'd0;
    mem[2828] = 'd1020;
    mem[2829] = 'd0;
    mem[2830] = 'd1020;
    mem[2831] = 'd0;
    mem[2832] = 'd0;
    mem[2833] = 'd0;
    mem[2834] = 'd1020;
    mem[2835] = 'd0;
    mem[2836] = 'd1020;
    mem[2837] = 'd0;
    mem[2838] = 'd0;
    mem[2839] = 'd0;
    mem[2840] = 'd912;
    mem[2841] = 'd0;
    mem[2842] = 'd964;
    mem[2843] = 'd0;
    mem[2844] = 'd0;
    mem[2845] = 'd0;
    mem[2846] = 'd188;
    mem[2847] = 'd0;
    mem[2848] = 'd648;
    mem[2849] = 'd0;
    mem[2850] = 'd0;
    mem[2851] = 'd0;
    mem[2852] = 'd32;
    mem[2853] = 'd0;
    mem[2854] = 'd708;
    mem[2855] = 'd0;
    mem[2856] = 'd0;
    mem[2857] = 'd0;
    mem[2858] = 'd220;
    mem[2859] = 'd0;
    mem[2860] = 'd836;
    mem[2861] = 'd0;
    mem[2862] = 'd0;
    mem[2863] = 'd0;
    mem[2864] = 'd632;
    mem[2865] = 'd0;
    mem[2866] = 'd976;
    mem[2867] = 'd0;
    mem[2868] = 'd0;
    mem[2869] = 'd0;
    mem[2870] = 'd696;
    mem[2871] = 'd0;
    mem[2872] = 'd1004;
    mem[2873] = 'd0;
    mem[2874] = 'd0;
    mem[2875] = 'd0;
    mem[2876] = 'd708;
    mem[2877] = 'd0;
    mem[2878] = 'd1004;
    mem[2879] = 'd0;
    mem[2880] = 'd0;
    mem[2881] = 'd0;
    mem[2882] = 'd720;
    mem[2883] = 'd0;
    mem[2884] = 'd1004;
    mem[2885] = 'd0;
    mem[2886] = 'd0;
    mem[2887] = 'd0;
    mem[2888] = 'd736;
    mem[2889] = 'd0;
    mem[2890] = 'd1004;
    mem[2891] = 'd0;
    mem[2892] = 'd0;
    mem[2893] = 'd0;
    mem[2894] = 'd752;
    mem[2895] = 'd0;
    mem[2896] = 'd1004;
    mem[2897] = 'd0;
    mem[2898] = 'd0;
    mem[2899] = 'd0;
    mem[2900] = 'd764;
    mem[2901] = 'd0;
    mem[2902] = 'd1004;
    mem[2903] = 'd0;
    mem[2904] = 'd0;
    mem[2905] = 'd0;
    mem[2906] = 'd780;
    mem[2907] = 'd0;
    mem[2908] = 'd1004;
    mem[2909] = 'd0;
    mem[2910] = 'd0;
    mem[2911] = 'd0;
    mem[2912] = 'd788;
    mem[2913] = 'd0;
    mem[2914] = 'd1008;
    mem[2915] = 'd0;
    mem[2916] = 'd0;
    mem[2917] = 'd0;
    mem[2918] = 'd796;
    mem[2919] = 'd0;
    mem[2920] = 'd1008;
    mem[2921] = 'd0;
    mem[2922] = 'd0;
    mem[2923] = 'd0;
    mem[2924] = 'd792;
    mem[2925] = 'd0;
    mem[2926] = 'd1008;
    mem[2927] = 'd0;
    mem[2928] = 'd0;
    mem[2929] = 'd0;
    mem[2930] = 'd788;
    mem[2931] = 'd0;
    mem[2932] = 'd1004;
    mem[2933] = 'd0;
    mem[2934] = 'd0;
    mem[2935] = 'd0;
    mem[2936] = 'd780;
    mem[2937] = 'd0;
    mem[2938] = 'd1004;
    mem[2939] = 'd0;
    mem[2940] = 'd0;
    mem[2941] = 'd0;
    mem[2942] = 'd764;
    mem[2943] = 'd0;
    mem[2944] = 'd1004;
    mem[2945] = 'd0;
    mem[2946] = 'd0;
    mem[2947] = 'd0;
    mem[2948] = 'd748;
    mem[2949] = 'd0;
    mem[2950] = 'd1004;
    mem[2951] = 'd0;
    mem[2952] = 'd0;
    mem[2953] = 'd0;
    mem[2954] = 'd732;
    mem[2955] = 'd0;
    mem[2956] = 'd1004;
    mem[2957] = 'd0;
    mem[2958] = 'd0;
    mem[2959] = 'd0;
    mem[2960] = 'd716;
    mem[2961] = 'd0;
    mem[2962] = 'd1004;
    mem[2963] = 'd0;
    mem[2964] = 'd0;
    mem[2965] = 'd0;
    mem[2966] = 'd704;
    mem[2967] = 'd0;
    mem[2968] = 'd1004;
    mem[2969] = 'd0;
    mem[2970] = 'd0;
    mem[2971] = 'd0;
    mem[2972] = 'd692;
    mem[2973] = 'd0;
    mem[2974] = 'd1004;
    mem[2975] = 'd0;
    mem[2976] = 'd0;
    mem[2977] = 'd0;
    mem[2978] = 'd656;
    mem[2979] = 'd0;
    mem[2980] = 'd980;
    mem[2981] = 'd0;
    mem[2982] = 'd0;
    mem[2983] = 'd0;
    mem[2984] = 'd300;
    mem[2985] = 'd0;
    mem[2986] = 'd860;
    mem[2987] = 'd0;
    mem[2988] = 'd0;
    mem[2989] = 'd0;
    mem[2990] = 'd32;
    mem[2991] = 'd0;
    mem[2992] = 'd708;
    mem[2993] = 'd0;
    mem[2994] = 'd0;
    mem[2995] = 'd0;
    mem[2996] = 'd160;
    mem[2997] = 'd0;
    mem[2998] = 'd644;
    mem[2999] = 'd0;
    mem[3000] = 'd0;
    mem[3001] = 'd0;
    mem[3002] = 'd904;
    mem[3003] = 'd0;
    mem[3004] = 'd960;
    mem[3005] = 'd0;
    mem[3006] = 'd0;
    mem[3007] = 'd0;
    mem[3008] = 'd1020;
    mem[3009] = 'd0;
    mem[3010] = 'd1020;
    mem[3011] = 'd0;
    mem[3012] = 'd0;
    mem[3013] = 'd0;
    mem[3014] = 'd1020;
    mem[3015] = 'd0;
    mem[3016] = 'd1020;
    mem[3017] = 'd0;
    mem[3018] = 'd0;
    mem[3019] = 'd0;
    mem[3020] = 'd1020;
    mem[3021] = 'd0;
    mem[3022] = 'd1020;
    mem[3023] = 'd0;
    mem[3024] = 'd0;
    mem[3025] = 'd0;
    mem[3026] = 'd1020;
    mem[3027] = 'd0;
    mem[3028] = 'd1020;
    mem[3029] = 'd0;
    mem[3030] = 'd0;
    mem[3031] = 'd0;
    mem[3032] = 'd1020;
    mem[3033] = 'd0;
    mem[3034] = 'd1020;
    mem[3035] = 'd0;
    mem[3036] = 'd0;
    mem[3037] = 'd0;
    mem[3038] = 'd1020;
    mem[3039] = 'd0;
    mem[3040] = 'd1020;
    mem[3041] = 'd0;
    mem[3042] = 'd0;
    mem[3043] = 'd1020;
    mem[3044] = 'd0;
    mem[3045] = 'd1020;
    mem[3046] = 'd0;
    mem[3047] = 'd0;
    mem[3048] = 'd0;
    mem[3049] = 'd1020;
    mem[3050] = 'd0;
    mem[3051] = 'd1020;
    mem[3052] = 'd0;
    mem[3053] = 'd0;
    mem[3054] = 'd0;
    mem[3055] = 'd1020;
    mem[3056] = 'd0;
    mem[3057] = 'd1020;
    mem[3058] = 'd0;
    mem[3059] = 'd0;
    mem[3060] = 'd0;
    mem[3061] = 'd1020;
    mem[3062] = 'd0;
    mem[3063] = 'd1020;
    mem[3064] = 'd0;
    mem[3065] = 'd0;
    mem[3066] = 'd0;
    mem[3067] = 'd1020;
    mem[3068] = 'd0;
    mem[3069] = 'd1020;
    mem[3070] = 'd0;
    mem[3071] = 'd0;
    mem[3072] = 'd0;
    mem[3073] = 'd964;
    mem[3074] = 'd0;
    mem[3075] = 'd1008;
    mem[3076] = 'd0;
    mem[3077] = 'd0;
    mem[3078] = 'd0;
    mem[3079] = 'd648;
    mem[3080] = 'd0;
    mem[3081] = 'd992;
    mem[3082] = 'd0;
    mem[3083] = 'd0;
    mem[3084] = 'd0;
    mem[3085] = 'd708;
    mem[3086] = 'd0;
    mem[3087] = 'd1020;
    mem[3088] = 'd0;
    mem[3089] = 'd0;
    mem[3090] = 'd0;
    mem[3091] = 'd836;
    mem[3092] = 'd0;
    mem[3093] = 'd1020;
    mem[3094] = 'd0;
    mem[3095] = 'd0;
    mem[3096] = 'd0;
    mem[3097] = 'd976;
    mem[3098] = 'd0;
    mem[3099] = 'd1020;
    mem[3100] = 'd0;
    mem[3101] = 'd0;
    mem[3102] = 'd0;
    mem[3103] = 'd1004;
    mem[3104] = 'd0;
    mem[3105] = 'd1020;
    mem[3106] = 'd0;
    mem[3107] = 'd0;
    mem[3108] = 'd0;
    mem[3109] = 'd1004;
    mem[3110] = 'd0;
    mem[3111] = 'd1020;
    mem[3112] = 'd0;
    mem[3113] = 'd0;
    mem[3114] = 'd0;
    mem[3115] = 'd1004;
    mem[3116] = 'd0;
    mem[3117] = 'd1020;
    mem[3118] = 'd0;
    mem[3119] = 'd0;
    mem[3120] = 'd0;
    mem[3121] = 'd1004;
    mem[3122] = 'd0;
    mem[3123] = 'd1020;
    mem[3124] = 'd0;
    mem[3125] = 'd0;
    mem[3126] = 'd0;
    mem[3127] = 'd1004;
    mem[3128] = 'd0;
    mem[3129] = 'd1020;
    mem[3130] = 'd0;
    mem[3131] = 'd0;
    mem[3132] = 'd0;
    mem[3133] = 'd1004;
    mem[3134] = 'd0;
    mem[3135] = 'd1020;
    mem[3136] = 'd0;
    mem[3137] = 'd0;
    mem[3138] = 'd0;
    mem[3139] = 'd1004;
    mem[3140] = 'd0;
    mem[3141] = 'd1020;
    mem[3142] = 'd0;
    mem[3143] = 'd0;
    mem[3144] = 'd0;
    mem[3145] = 'd1008;
    mem[3146] = 'd0;
    mem[3147] = 'd1020;
    mem[3148] = 'd0;
    mem[3149] = 'd0;
    mem[3150] = 'd0;
    mem[3151] = 'd1008;
    mem[3152] = 'd0;
    mem[3153] = 'd1020;
    mem[3154] = 'd0;
    mem[3155] = 'd0;
    mem[3156] = 'd0;
    mem[3157] = 'd1008;
    mem[3158] = 'd0;
    mem[3159] = 'd1020;
    mem[3160] = 'd0;
    mem[3161] = 'd0;
    mem[3162] = 'd0;
    mem[3163] = 'd1004;
    mem[3164] = 'd0;
    mem[3165] = 'd1020;
    mem[3166] = 'd0;
    mem[3167] = 'd0;
    mem[3168] = 'd0;
    mem[3169] = 'd1004;
    mem[3170] = 'd0;
    mem[3171] = 'd1020;
    mem[3172] = 'd0;
    mem[3173] = 'd0;
    mem[3174] = 'd0;
    mem[3175] = 'd1004;
    mem[3176] = 'd0;
    mem[3177] = 'd1020;
    mem[3178] = 'd0;
    mem[3179] = 'd0;
    mem[3180] = 'd0;
    mem[3181] = 'd1004;
    mem[3182] = 'd0;
    mem[3183] = 'd1020;
    mem[3184] = 'd0;
    mem[3185] = 'd0;
    mem[3186] = 'd0;
    mem[3187] = 'd1004;
    mem[3188] = 'd0;
    mem[3189] = 'd1020;
    mem[3190] = 'd0;
    mem[3191] = 'd0;
    mem[3192] = 'd0;
    mem[3193] = 'd1004;
    mem[3194] = 'd0;
    mem[3195] = 'd1020;
    mem[3196] = 'd0;
    mem[3197] = 'd0;
    mem[3198] = 'd0;
    mem[3199] = 'd1004;
    mem[3200] = 'd0;
    mem[3201] = 'd1020;
    mem[3202] = 'd0;
    mem[3203] = 'd0;
    mem[3204] = 'd0;
    mem[3205] = 'd1004;
    mem[3206] = 'd0;
    mem[3207] = 'd1020;
    mem[3208] = 'd0;
    mem[3209] = 'd0;
    mem[3210] = 'd0;
    mem[3211] = 'd980;
    mem[3212] = 'd0;
    mem[3213] = 'd1020;
    mem[3214] = 'd0;
    mem[3215] = 'd0;
    mem[3216] = 'd0;
    mem[3217] = 'd860;
    mem[3218] = 'd0;
    mem[3219] = 'd1020;
    mem[3220] = 'd0;
    mem[3221] = 'd0;
    mem[3222] = 'd0;
    mem[3223] = 'd708;
    mem[3224] = 'd0;
    mem[3225] = 'd1020;
    mem[3226] = 'd0;
    mem[3227] = 'd0;
    mem[3228] = 'd0;
    mem[3229] = 'd644;
    mem[3230] = 'd0;
    mem[3231] = 'd996;
    mem[3232] = 'd0;
    mem[3233] = 'd0;
    mem[3234] = 'd0;
    mem[3235] = 'd960;
    mem[3236] = 'd0;
    mem[3237] = 'd1012;
    mem[3238] = 'd0;
    mem[3239] = 'd0;
    mem[3240] = 'd0;
    mem[3241] = 'd1020;
    mem[3242] = 'd0;
    mem[3243] = 'd1020;
    mem[3244] = 'd0;
    mem[3245] = 'd0;
    mem[3246] = 'd0;
    mem[3247] = 'd1020;
    mem[3248] = 'd0;
    mem[3249] = 'd1020;
    mem[3250] = 'd0;
    mem[3251] = 'd0;
    mem[3252] = 'd0;
    mem[3253] = 'd1020;
    mem[3254] = 'd0;
    mem[3255] = 'd1020;
    mem[3256] = 'd0;
    mem[3257] = 'd0;
    mem[3258] = 'd0;
    mem[3259] = 'd1020;
    mem[3260] = 'd0;
    mem[3261] = 'd1020;
    mem[3262] = 'd0;
    mem[3263] = 'd0;
    mem[3264] = 'd0;
    mem[3265] = 'd1020;
    mem[3266] = 'd0;
    mem[3267] = 'd1020;
    mem[3268] = 'd0;
    mem[3269] = 'd0;
    mem[3270] = 'd0;
    mem[3271] = 'd1020;
    mem[3272] = 'd0;
    mem[3273] = 'd1020;
    mem[3274] = 'd0;
    mem[3275] = 'd0;
    mem[3276] = 'd0;
    mem[3277] = 'd0;
    mem[3278] = 'd1020;
    mem[3279] = 'd0;
    mem[3280] = 'd1020;
    mem[3281] = 'd0;
    mem[3282] = 'd0;
    mem[3283] = 'd0;
    mem[3284] = 'd1020;
    mem[3285] = 'd0;
    mem[3286] = 'd1020;
    mem[3287] = 'd0;
    mem[3288] = 'd0;
    mem[3289] = 'd0;
    mem[3290] = 'd1020;
    mem[3291] = 'd0;
    mem[3292] = 'd1020;
    mem[3293] = 'd0;
    mem[3294] = 'd0;
    mem[3295] = 'd0;
    mem[3296] = 'd1020;
    mem[3297] = 'd0;
    mem[3298] = 'd1020;
    mem[3299] = 'd0;
    mem[3300] = 'd0;
    mem[3301] = 'd0;
    mem[3302] = 'd964;
    mem[3303] = 'd0;
    mem[3304] = 'd984;
    mem[3305] = 'd0;
    mem[3306] = 'd0;
    mem[3307] = 'd0;
    mem[3308] = 'd248;
    mem[3309] = 'd0;
    mem[3310] = 'd660;
    mem[3311] = 'd0;
    mem[3312] = 'd0;
    mem[3313] = 'd0;
    mem[3314] = 'd32;
    mem[3315] = 'd0;
    mem[3316] = 'd688;
    mem[3317] = 'd0;
    mem[3318] = 'd0;
    mem[3319] = 'd0;
    mem[3320] = 'd232;
    mem[3321] = 'd0;
    mem[3322] = 'd832;
    mem[3323] = 'd0;
    mem[3324] = 'd0;
    mem[3325] = 'd0;
    mem[3326] = 'd592;
    mem[3327] = 'd0;
    mem[3328] = 'd960;
    mem[3329] = 'd0;
    mem[3330] = 'd0;
    mem[3331] = 'd0;
    mem[3332] = 'd628;
    mem[3333] = 'd0;
    mem[3334] = 'd988;
    mem[3335] = 'd0;
    mem[3336] = 'd0;
    mem[3337] = 'd0;
    mem[3338] = 'd640;
    mem[3339] = 'd0;
    mem[3340] = 'd996;
    mem[3341] = 'd0;
    mem[3342] = 'd0;
    mem[3343] = 'd0;
    mem[3344] = 'd652;
    mem[3345] = 'd0;
    mem[3346] = 'd1000;
    mem[3347] = 'd0;
    mem[3348] = 'd0;
    mem[3349] = 'd0;
    mem[3350] = 'd664;
    mem[3351] = 'd0;
    mem[3352] = 'd1000;
    mem[3353] = 'd0;
    mem[3354] = 'd0;
    mem[3355] = 'd0;
    mem[3356] = 'd676;
    mem[3357] = 'd0;
    mem[3358] = 'd1000;
    mem[3359] = 'd0;
    mem[3360] = 'd0;
    mem[3361] = 'd0;
    mem[3362] = 'd692;
    mem[3363] = 'd0;
    mem[3364] = 'd1004;
    mem[3365] = 'd0;
    mem[3366] = 'd0;
    mem[3367] = 'd0;
    mem[3368] = 'd708;
    mem[3369] = 'd0;
    mem[3370] = 'd1004;
    mem[3371] = 'd0;
    mem[3372] = 'd0;
    mem[3373] = 'd0;
    mem[3374] = 'd716;
    mem[3375] = 'd0;
    mem[3376] = 'd1004;
    mem[3377] = 'd0;
    mem[3378] = 'd0;
    mem[3379] = 'd0;
    mem[3380] = 'd728;
    mem[3381] = 'd0;
    mem[3382] = 'd1004;
    mem[3383] = 'd0;
    mem[3384] = 'd0;
    mem[3385] = 'd0;
    mem[3386] = 'd732;
    mem[3387] = 'd0;
    mem[3388] = 'd1004;
    mem[3389] = 'd0;
    mem[3390] = 'd0;
    mem[3391] = 'd0;
    mem[3392] = 'd732;
    mem[3393] = 'd0;
    mem[3394] = 'd1004;
    mem[3395] = 'd0;
    mem[3396] = 'd0;
    mem[3397] = 'd0;
    mem[3398] = 'd724;
    mem[3399] = 'd0;
    mem[3400] = 'd1004;
    mem[3401] = 'd0;
    mem[3402] = 'd0;
    mem[3403] = 'd0;
    mem[3404] = 'd716;
    mem[3405] = 'd0;
    mem[3406] = 'd1004;
    mem[3407] = 'd0;
    mem[3408] = 'd0;
    mem[3409] = 'd0;
    mem[3410] = 'd704;
    mem[3411] = 'd0;
    mem[3412] = 'd1004;
    mem[3413] = 'd0;
    mem[3414] = 'd0;
    mem[3415] = 'd0;
    mem[3416] = 'd692;
    mem[3417] = 'd0;
    mem[3418] = 'd1004;
    mem[3419] = 'd0;
    mem[3420] = 'd0;
    mem[3421] = 'd0;
    mem[3422] = 'd676;
    mem[3423] = 'd0;
    mem[3424] = 'd1000;
    mem[3425] = 'd0;
    mem[3426] = 'd0;
    mem[3427] = 'd0;
    mem[3428] = 'd664;
    mem[3429] = 'd0;
    mem[3430] = 'd1000;
    mem[3431] = 'd0;
    mem[3432] = 'd0;
    mem[3433] = 'd0;
    mem[3434] = 'd652;
    mem[3435] = 'd0;
    mem[3436] = 'd1000;
    mem[3437] = 'd0;
    mem[3438] = 'd0;
    mem[3439] = 'd0;
    mem[3440] = 'd640;
    mem[3441] = 'd0;
    mem[3442] = 'd996;
    mem[3443] = 'd0;
    mem[3444] = 'd0;
    mem[3445] = 'd0;
    mem[3446] = 'd628;
    mem[3447] = 'd0;
    mem[3448] = 'd988;
    mem[3449] = 'd0;
    mem[3450] = 'd0;
    mem[3451] = 'd0;
    mem[3452] = 'd616;
    mem[3453] = 'd0;
    mem[3454] = 'd964;
    mem[3455] = 'd0;
    mem[3456] = 'd0;
    mem[3457] = 'd0;
    mem[3458] = 'd300;
    mem[3459] = 'd0;
    mem[3460] = 'd852;
    mem[3461] = 'd0;
    mem[3462] = 'd0;
    mem[3463] = 'd0;
    mem[3464] = 'd28;
    mem[3465] = 'd0;
    mem[3466] = 'd692;
    mem[3467] = 'd0;
    mem[3468] = 'd0;
    mem[3469] = 'd0;
    mem[3470] = 'd212;
    mem[3471] = 'd0;
    mem[3472] = 'd648;
    mem[3473] = 'd0;
    mem[3474] = 'd0;
    mem[3475] = 'd0;
    mem[3476] = 'd948;
    mem[3477] = 'd0;
    mem[3478] = 'd976;
    mem[3479] = 'd0;
    mem[3480] = 'd0;
    mem[3481] = 'd0;
    mem[3482] = 'd1020;
    mem[3483] = 'd0;
    mem[3484] = 'd1020;
    mem[3485] = 'd0;
    mem[3486] = 'd0;
    mem[3487] = 'd0;
    mem[3488] = 'd1020;
    mem[3489] = 'd0;
    mem[3490] = 'd1020;
    mem[3491] = 'd0;
    mem[3492] = 'd0;
    mem[3493] = 'd0;
    mem[3494] = 'd1020;
    mem[3495] = 'd0;
    mem[3496] = 'd1020;
    mem[3497] = 'd0;
    mem[3498] = 'd0;
    mem[3499] = 'd0;
    mem[3500] = 'd1020;
    mem[3501] = 'd0;
    mem[3502] = 'd1020;
    mem[3503] = 'd0;
    mem[3504] = 'd0;
    mem[3505] = 'd0;
    mem[3506] = 'd1020;
    mem[3507] = 'd0;
    mem[3508] = 'd1020;
    mem[3509] = 'd0;
    mem[3510] = 'd0;
    mem[3511] = 'd1020;
    mem[3512] = 'd0;
    mem[3513] = 'd1020;
    mem[3514] = 'd0;
    mem[3515] = 'd0;
    mem[3516] = 'd0;
    mem[3517] = 'd1020;
    mem[3518] = 'd0;
    mem[3519] = 'd1020;
    mem[3520] = 'd0;
    mem[3521] = 'd0;
    mem[3522] = 'd0;
    mem[3523] = 'd1020;
    mem[3524] = 'd0;
    mem[3525] = 'd1020;
    mem[3526] = 'd0;
    mem[3527] = 'd0;
    mem[3528] = 'd0;
    mem[3529] = 'd1020;
    mem[3530] = 'd0;
    mem[3531] = 'd1020;
    mem[3532] = 'd0;
    mem[3533] = 'd0;
    mem[3534] = 'd0;
    mem[3535] = 'd984;
    mem[3536] = 'd0;
    mem[3537] = 'd1004;
    mem[3538] = 'd0;
    mem[3539] = 'd0;
    mem[3540] = 'd0;
    mem[3541] = 'd660;
    mem[3542] = 'd0;
    mem[3543] = 'd980;
    mem[3544] = 'd0;
    mem[3545] = 'd0;
    mem[3546] = 'd0;
    mem[3547] = 'd688;
    mem[3548] = 'd0;
    mem[3549] = 'd1020;
    mem[3550] = 'd0;
    mem[3551] = 'd0;
    mem[3552] = 'd0;
    mem[3553] = 'd832;
    mem[3554] = 'd0;
    mem[3555] = 'd1020;
    mem[3556] = 'd0;
    mem[3557] = 'd0;
    mem[3558] = 'd0;
    mem[3559] = 'd960;
    mem[3560] = 'd0;
    mem[3561] = 'd1020;
    mem[3562] = 'd0;
    mem[3563] = 'd0;
    mem[3564] = 'd0;
    mem[3565] = 'd988;
    mem[3566] = 'd0;
    mem[3567] = 'd1020;
    mem[3568] = 'd0;
    mem[3569] = 'd0;
    mem[3570] = 'd0;
    mem[3571] = 'd996;
    mem[3572] = 'd0;
    mem[3573] = 'd1020;
    mem[3574] = 'd0;
    mem[3575] = 'd0;
    mem[3576] = 'd0;
    mem[3577] = 'd1000;
    mem[3578] = 'd0;
    mem[3579] = 'd1020;
    mem[3580] = 'd0;
    mem[3581] = 'd0;
    mem[3582] = 'd0;
    mem[3583] = 'd1000;
    mem[3584] = 'd0;
    mem[3585] = 'd1020;
    mem[3586] = 'd0;
    mem[3587] = 'd0;
    mem[3588] = 'd0;
    mem[3589] = 'd1000;
    mem[3590] = 'd0;
    mem[3591] = 'd1020;
    mem[3592] = 'd0;
    mem[3593] = 'd0;
    mem[3594] = 'd0;
    mem[3595] = 'd1004;
    mem[3596] = 'd0;
    mem[3597] = 'd1020;
    mem[3598] = 'd0;
    mem[3599] = 'd0;
    mem[3600] = 'd0;
    mem[3601] = 'd1004;
    mem[3602] = 'd0;
    mem[3603] = 'd1020;
    mem[3604] = 'd0;
    mem[3605] = 'd0;
    mem[3606] = 'd0;
    mem[3607] = 'd1004;
    mem[3608] = 'd0;
    mem[3609] = 'd1020;
    mem[3610] = 'd0;
    mem[3611] = 'd0;
    mem[3612] = 'd0;
    mem[3613] = 'd1004;
    mem[3614] = 'd0;
    mem[3615] = 'd1020;
    mem[3616] = 'd0;
    mem[3617] = 'd0;
    mem[3618] = 'd0;
    mem[3619] = 'd1004;
    mem[3620] = 'd0;
    mem[3621] = 'd1020;
    mem[3622] = 'd0;
    mem[3623] = 'd0;
    mem[3624] = 'd0;
    mem[3625] = 'd1004;
    mem[3626] = 'd0;
    mem[3627] = 'd1020;
    mem[3628] = 'd0;
    mem[3629] = 'd0;
    mem[3630] = 'd0;
    mem[3631] = 'd1004;
    mem[3632] = 'd0;
    mem[3633] = 'd1020;
    mem[3634] = 'd0;
    mem[3635] = 'd0;
    mem[3636] = 'd0;
    mem[3637] = 'd1004;
    mem[3638] = 'd0;
    mem[3639] = 'd1020;
    mem[3640] = 'd0;
    mem[3641] = 'd0;
    mem[3642] = 'd0;
    mem[3643] = 'd1004;
    mem[3644] = 'd0;
    mem[3645] = 'd1020;
    mem[3646] = 'd0;
    mem[3647] = 'd0;
    mem[3648] = 'd0;
    mem[3649] = 'd1004;
    mem[3650] = 'd0;
    mem[3651] = 'd1020;
    mem[3652] = 'd0;
    mem[3653] = 'd0;
    mem[3654] = 'd0;
    mem[3655] = 'd1000;
    mem[3656] = 'd0;
    mem[3657] = 'd1020;
    mem[3658] = 'd0;
    mem[3659] = 'd0;
    mem[3660] = 'd0;
    mem[3661] = 'd1000;
    mem[3662] = 'd0;
    mem[3663] = 'd1020;
    mem[3664] = 'd0;
    mem[3665] = 'd0;
    mem[3666] = 'd0;
    mem[3667] = 'd1000;
    mem[3668] = 'd0;
    mem[3669] = 'd1020;
    mem[3670] = 'd0;
    mem[3671] = 'd0;
    mem[3672] = 'd0;
    mem[3673] = 'd996;
    mem[3674] = 'd0;
    mem[3675] = 'd1020;
    mem[3676] = 'd0;
    mem[3677] = 'd0;
    mem[3678] = 'd0;
    mem[3679] = 'd988;
    mem[3680] = 'd0;
    mem[3681] = 'd1020;
    mem[3682] = 'd0;
    mem[3683] = 'd0;
    mem[3684] = 'd0;
    mem[3685] = 'd964;
    mem[3686] = 'd0;
    mem[3687] = 'd1020;
    mem[3688] = 'd0;
    mem[3689] = 'd0;
    mem[3690] = 'd0;
    mem[3691] = 'd852;
    mem[3692] = 'd0;
    mem[3693] = 'd1020;
    mem[3694] = 'd0;
    mem[3695] = 'd0;
    mem[3696] = 'd0;
    mem[3697] = 'd692;
    mem[3698] = 'd0;
    mem[3699] = 'd1020;
    mem[3700] = 'd0;
    mem[3701] = 'd0;
    mem[3702] = 'd0;
    mem[3703] = 'd648;
    mem[3704] = 'd0;
    mem[3705] = 'd984;
    mem[3706] = 'd0;
    mem[3707] = 'd0;
    mem[3708] = 'd0;
    mem[3709] = 'd976;
    mem[3710] = 'd0;
    mem[3711] = 'd1004;
    mem[3712] = 'd0;
    mem[3713] = 'd0;
    mem[3714] = 'd0;
    mem[3715] = 'd1020;
    mem[3716] = 'd0;
    mem[3717] = 'd1020;
    mem[3718] = 'd0;
    mem[3719] = 'd0;
    mem[3720] = 'd0;
    mem[3721] = 'd1020;
    mem[3722] = 'd0;
    mem[3723] = 'd1020;
    mem[3724] = 'd0;
    mem[3725] = 'd0;
    mem[3726] = 'd0;
    mem[3727] = 'd1020;
    mem[3728] = 'd0;
    mem[3729] = 'd1020;
    mem[3730] = 'd0;
    mem[3731] = 'd0;
    mem[3732] = 'd0;
    mem[3733] = 'd1020;
    mem[3734] = 'd0;
    mem[3735] = 'd1020;
    mem[3736] = 'd0;
    mem[3737] = 'd0;
    mem[3738] = 'd0;
    mem[3739] = 'd1020;
    mem[3740] = 'd0;
    mem[3741] = 'd1020;
    mem[3742] = 'd0;
    mem[3743] = 'd0;
    mem[3744] = 'd0;
    mem[3745] = 'd0;
    mem[3746] = 'd1020;
    mem[3747] = 'd0;
    mem[3748] = 'd1020;
    mem[3749] = 'd0;
    mem[3750] = 'd0;
    mem[3751] = 'd0;
    mem[3752] = 'd1020;
    mem[3753] = 'd0;
    mem[3754] = 'd1020;
    mem[3755] = 'd0;
    mem[3756] = 'd0;
    mem[3757] = 'd0;
    mem[3758] = 'd1020;
    mem[3759] = 'd0;
    mem[3760] = 'd1020;
    mem[3761] = 'd0;
    mem[3762] = 'd0;
    mem[3763] = 'd0;
    mem[3764] = 'd1020;
    mem[3765] = 'd0;
    mem[3766] = 'd1020;
    mem[3767] = 'd0;
    mem[3768] = 'd0;
    mem[3769] = 'd0;
    mem[3770] = 'd452;
    mem[3771] = 'd0;
    mem[3772] = 'd748;
    mem[3773] = 'd0;
    mem[3774] = 'd0;
    mem[3775] = 'd0;
    mem[3776] = 'd24;
    mem[3777] = 'd0;
    mem[3778] = 'd656;
    mem[3779] = 'd0;
    mem[3780] = 'd0;
    mem[3781] = 'd0;
    mem[3782] = 'd160;
    mem[3783] = 'd0;
    mem[3784] = 'd796;
    mem[3785] = 'd0;
    mem[3786] = 'd0;
    mem[3787] = 'd0;
    mem[3788] = 'd524;
    mem[3789] = 'd0;
    mem[3790] = 'd932;
    mem[3791] = 'd0;
    mem[3792] = 'd0;
    mem[3793] = 'd0;
    mem[3794] = 'd560;
    mem[3795] = 'd0;
    mem[3796] = 'd964;
    mem[3797] = 'd0;
    mem[3798] = 'd0;
    mem[3799] = 'd0;
    mem[3800] = 'd572;
    mem[3801] = 'd0;
    mem[3802] = 'd984;
    mem[3803] = 'd0;
    mem[3804] = 'd0;
    mem[3805] = 'd0;
    mem[3806] = 'd584;
    mem[3807] = 'd0;
    mem[3808] = 'd996;
    mem[3809] = 'd0;
    mem[3810] = 'd0;
    mem[3811] = 'd0;
    mem[3812] = 'd592;
    mem[3813] = 'd0;
    mem[3814] = 'd996;
    mem[3815] = 'd0;
    mem[3816] = 'd0;
    mem[3817] = 'd0;
    mem[3818] = 'd604;
    mem[3819] = 'd0;
    mem[3820] = 'd996;
    mem[3821] = 'd0;
    mem[3822] = 'd0;
    mem[3823] = 'd0;
    mem[3824] = 'd616;
    mem[3825] = 'd0;
    mem[3826] = 'd996;
    mem[3827] = 'd0;
    mem[3828] = 'd0;
    mem[3829] = 'd0;
    mem[3830] = 'd628;
    mem[3831] = 'd0;
    mem[3832] = 'd996;
    mem[3833] = 'd0;
    mem[3834] = 'd0;
    mem[3835] = 'd0;
    mem[3836] = 'd644;
    mem[3837] = 'd0;
    mem[3838] = 'd1000;
    mem[3839] = 'd0;
    mem[3840] = 'd0;
    mem[3841] = 'd0;
    mem[3842] = 'd652;
    mem[3843] = 'd0;
    mem[3844] = 'd1000;
    mem[3845] = 'd0;
    mem[3846] = 'd0;
    mem[3847] = 'd0;
    mem[3848] = 'd660;
    mem[3849] = 'd0;
    mem[3850] = 'd1000;
    mem[3851] = 'd0;
    mem[3852] = 'd0;
    mem[3853] = 'd0;
    mem[3854] = 'd664;
    mem[3855] = 'd0;
    mem[3856] = 'd1000;
    mem[3857] = 'd0;
    mem[3858] = 'd0;
    mem[3859] = 'd0;
    mem[3860] = 'd664;
    mem[3861] = 'd0;
    mem[3862] = 'd1000;
    mem[3863] = 'd0;
    mem[3864] = 'd0;
    mem[3865] = 'd0;
    mem[3866] = 'd660;
    mem[3867] = 'd0;
    mem[3868] = 'd1000;
    mem[3869] = 'd0;
    mem[3870] = 'd0;
    mem[3871] = 'd0;
    mem[3872] = 'd652;
    mem[3873] = 'd0;
    mem[3874] = 'd1000;
    mem[3875] = 'd0;
    mem[3876] = 'd0;
    mem[3877] = 'd0;
    mem[3878] = 'd640;
    mem[3879] = 'd0;
    mem[3880] = 'd1000;
    mem[3881] = 'd0;
    mem[3882] = 'd0;
    mem[3883] = 'd0;
    mem[3884] = 'd628;
    mem[3885] = 'd0;
    mem[3886] = 'd996;
    mem[3887] = 'd0;
    mem[3888] = 'd0;
    mem[3889] = 'd0;
    mem[3890] = 'd616;
    mem[3891] = 'd0;
    mem[3892] = 'd996;
    mem[3893] = 'd0;
    mem[3894] = 'd0;
    mem[3895] = 'd0;
    mem[3896] = 'd604;
    mem[3897] = 'd0;
    mem[3898] = 'd996;
    mem[3899] = 'd0;
    mem[3900] = 'd0;
    mem[3901] = 'd0;
    mem[3902] = 'd592;
    mem[3903] = 'd0;
    mem[3904] = 'd996;
    mem[3905] = 'd0;
    mem[3906] = 'd0;
    mem[3907] = 'd0;
    mem[3908] = 'd584;
    mem[3909] = 'd0;
    mem[3910] = 'd996;
    mem[3911] = 'd0;
    mem[3912] = 'd0;
    mem[3913] = 'd0;
    mem[3914] = 'd572;
    mem[3915] = 'd0;
    mem[3916] = 'd988;
    mem[3917] = 'd0;
    mem[3918] = 'd0;
    mem[3919] = 'd0;
    mem[3920] = 'd560;
    mem[3921] = 'd0;
    mem[3922] = 'd968;
    mem[3923] = 'd0;
    mem[3924] = 'd0;
    mem[3925] = 'd0;
    mem[3926] = 'd544;
    mem[3927] = 'd0;
    mem[3928] = 'd936;
    mem[3929] = 'd0;
    mem[3930] = 'd0;
    mem[3931] = 'd0;
    mem[3932] = 'd232;
    mem[3933] = 'd0;
    mem[3934] = 'd812;
    mem[3935] = 'd0;
    mem[3936] = 'd0;
    mem[3937] = 'd0;
    mem[3938] = 'd24;
    mem[3939] = 'd0;
    mem[3940] = 'd660;
    mem[3941] = 'd0;
    mem[3942] = 'd0;
    mem[3943] = 'd0;
    mem[3944] = 'd468;
    mem[3945] = 'd0;
    mem[3946] = 'd752;
    mem[3947] = 'd0;
    mem[3948] = 'd0;
    mem[3949] = 'd0;
    mem[3950] = 'd1020;
    mem[3951] = 'd0;
    mem[3952] = 'd1020;
    mem[3953] = 'd0;
    mem[3954] = 'd0;
    mem[3955] = 'd0;
    mem[3956] = 'd1020;
    mem[3957] = 'd0;
    mem[3958] = 'd1020;
    mem[3959] = 'd0;
    mem[3960] = 'd0;
    mem[3961] = 'd0;
    mem[3962] = 'd1020;
    mem[3963] = 'd0;
    mem[3964] = 'd1020;
    mem[3965] = 'd0;
    mem[3966] = 'd0;
    mem[3967] = 'd0;
    mem[3968] = 'd1020;
    mem[3969] = 'd0;
    mem[3970] = 'd1020;
    mem[3971] = 'd0;
    mem[3972] = 'd0;
    mem[3973] = 'd0;
    mem[3974] = 'd1020;
    mem[3975] = 'd0;
    mem[3976] = 'd1020;
    mem[3977] = 'd0;
    mem[3978] = 'd0;
    mem[3979] = 'd1020;
    mem[3980] = 'd0;
    mem[3981] = 'd1020;
    mem[3982] = 'd0;
    mem[3983] = 'd0;
    mem[3984] = 'd0;
    mem[3985] = 'd1020;
    mem[3986] = 'd0;
    mem[3987] = 'd1020;
    mem[3988] = 'd0;
    mem[3989] = 'd0;
    mem[3990] = 'd0;
    mem[3991] = 'd1020;
    mem[3992] = 'd0;
    mem[3993] = 'd1020;
    mem[3994] = 'd0;
    mem[3995] = 'd0;
    mem[3996] = 'd0;
    mem[3997] = 'd1020;
    mem[3998] = 'd0;
    mem[3999] = 'd1020;
    mem[4000] = 'd0;
    mem[4001] = 'd0;
    mem[4002] = 'd0;
    mem[4003] = 'd748;
    mem[4004] = 'd0;
    mem[4005] = 'd988;
    mem[4006] = 'd0;
    mem[4007] = 'd0;
    mem[4008] = 'd0;
    mem[4009] = 'd656;
    mem[4010] = 'd0;
    mem[4011] = 'd1020;
    mem[4012] = 'd0;
    mem[4013] = 'd0;
    mem[4014] = 'd0;
    mem[4015] = 'd796;
    mem[4016] = 'd0;
    mem[4017] = 'd1020;
    mem[4018] = 'd0;
    mem[4019] = 'd0;
    mem[4020] = 'd0;
    mem[4021] = 'd932;
    mem[4022] = 'd0;
    mem[4023] = 'd1020;
    mem[4024] = 'd0;
    mem[4025] = 'd0;
    mem[4026] = 'd0;
    mem[4027] = 'd964;
    mem[4028] = 'd0;
    mem[4029] = 'd1020;
    mem[4030] = 'd0;
    mem[4031] = 'd0;
    mem[4032] = 'd0;
    mem[4033] = 'd984;
    mem[4034] = 'd0;
    mem[4035] = 'd1020;
    mem[4036] = 'd0;
    mem[4037] = 'd0;
    mem[4038] = 'd0;
    mem[4039] = 'd996;
    mem[4040] = 'd0;
    mem[4041] = 'd1020;
    mem[4042] = 'd0;
    mem[4043] = 'd0;
    mem[4044] = 'd0;
    mem[4045] = 'd996;
    mem[4046] = 'd0;
    mem[4047] = 'd1020;
    mem[4048] = 'd0;
    mem[4049] = 'd0;
    mem[4050] = 'd0;
    mem[4051] = 'd996;
    mem[4052] = 'd0;
    mem[4053] = 'd1020;
    mem[4054] = 'd0;
    mem[4055] = 'd0;
    mem[4056] = 'd0;
    mem[4057] = 'd996;
    mem[4058] = 'd0;
    mem[4059] = 'd1020;
    mem[4060] = 'd0;
    mem[4061] = 'd0;
    mem[4062] = 'd0;
    mem[4063] = 'd996;
    mem[4064] = 'd0;
    mem[4065] = 'd1020;
    mem[4066] = 'd0;
    mem[4067] = 'd0;
    mem[4068] = 'd0;
    mem[4069] = 'd1000;
    mem[4070] = 'd0;
    mem[4071] = 'd1020;
    mem[4072] = 'd0;
    mem[4073] = 'd0;
    mem[4074] = 'd0;
    mem[4075] = 'd1000;
    mem[4076] = 'd0;
    mem[4077] = 'd1020;
    mem[4078] = 'd0;
    mem[4079] = 'd0;
    mem[4080] = 'd0;
    mem[4081] = 'd1000;
    mem[4082] = 'd0;
    mem[4083] = 'd1020;
    mem[4084] = 'd0;
    mem[4085] = 'd0;
    mem[4086] = 'd0;
    mem[4087] = 'd1000;
    mem[4088] = 'd0;
    mem[4089] = 'd1020;
    mem[4090] = 'd0;
    mem[4091] = 'd0;
    mem[4092] = 'd0;
    mem[4093] = 'd1000;
    mem[4094] = 'd0;
    mem[4095] = 'd1020;
    mem[4096] = 'd0;
    mem[4097] = 'd0;
    mem[4098] = 'd0;
    mem[4099] = 'd1000;
    mem[4100] = 'd0;
    mem[4101] = 'd1020;
    mem[4102] = 'd0;
    mem[4103] = 'd0;
    mem[4104] = 'd0;
    mem[4105] = 'd1000;
    mem[4106] = 'd0;
    mem[4107] = 'd1020;
    mem[4108] = 'd0;
    mem[4109] = 'd0;
    mem[4110] = 'd0;
    mem[4111] = 'd1000;
    mem[4112] = 'd0;
    mem[4113] = 'd1020;
    mem[4114] = 'd0;
    mem[4115] = 'd0;
    mem[4116] = 'd0;
    mem[4117] = 'd996;
    mem[4118] = 'd0;
    mem[4119] = 'd1020;
    mem[4120] = 'd0;
    mem[4121] = 'd0;
    mem[4122] = 'd0;
    mem[4123] = 'd996;
    mem[4124] = 'd0;
    mem[4125] = 'd1020;
    mem[4126] = 'd0;
    mem[4127] = 'd0;
    mem[4128] = 'd0;
    mem[4129] = 'd996;
    mem[4130] = 'd0;
    mem[4131] = 'd1020;
    mem[4132] = 'd0;
    mem[4133] = 'd0;
    mem[4134] = 'd0;
    mem[4135] = 'd996;
    mem[4136] = 'd0;
    mem[4137] = 'd1020;
    mem[4138] = 'd0;
    mem[4139] = 'd0;
    mem[4140] = 'd0;
    mem[4141] = 'd996;
    mem[4142] = 'd0;
    mem[4143] = 'd1020;
    mem[4144] = 'd0;
    mem[4145] = 'd0;
    mem[4146] = 'd0;
    mem[4147] = 'd988;
    mem[4148] = 'd0;
    mem[4149] = 'd1020;
    mem[4150] = 'd0;
    mem[4151] = 'd0;
    mem[4152] = 'd0;
    mem[4153] = 'd968;
    mem[4154] = 'd0;
    mem[4155] = 'd1020;
    mem[4156] = 'd0;
    mem[4157] = 'd0;
    mem[4158] = 'd0;
    mem[4159] = 'd936;
    mem[4160] = 'd0;
    mem[4161] = 'd1020;
    mem[4162] = 'd0;
    mem[4163] = 'd0;
    mem[4164] = 'd0;
    mem[4165] = 'd812;
    mem[4166] = 'd0;
    mem[4167] = 'd1020;
    mem[4168] = 'd0;
    mem[4169] = 'd0;
    mem[4170] = 'd0;
    mem[4171] = 'd660;
    mem[4172] = 'd0;
    mem[4173] = 'd1020;
    mem[4174] = 'd0;
    mem[4175] = 'd0;
    mem[4176] = 'd0;
    mem[4177] = 'd752;
    mem[4178] = 'd0;
    mem[4179] = 'd984;
    mem[4180] = 'd0;
    mem[4181] = 'd0;
    mem[4182] = 'd0;
    mem[4183] = 'd1020;
    mem[4184] = 'd0;
    mem[4185] = 'd1020;
    mem[4186] = 'd0;
    mem[4187] = 'd0;
    mem[4188] = 'd0;
    mem[4189] = 'd1020;
    mem[4190] = 'd0;
    mem[4191] = 'd1020;
    mem[4192] = 'd0;
    mem[4193] = 'd0;
    mem[4194] = 'd0;
    mem[4195] = 'd1020;
    mem[4196] = 'd0;
    mem[4197] = 'd1020;
    mem[4198] = 'd0;
    mem[4199] = 'd0;
    mem[4200] = 'd0;
    mem[4201] = 'd1020;
    mem[4202] = 'd0;
    mem[4203] = 'd1020;
    mem[4204] = 'd0;
    mem[4205] = 'd0;
    mem[4206] = 'd0;
    mem[4207] = 'd1020;
    mem[4208] = 'd0;
    mem[4209] = 'd1020;
    mem[4210] = 'd0;
    mem[4211] = 'd0;
    mem[4212] = 'd0;
    mem[4213] = 'd0;
    mem[4214] = 'd1020;
    mem[4215] = 'd0;
    mem[4216] = 'd1020;
    mem[4217] = 'd0;
    mem[4218] = 'd0;
    mem[4219] = 'd0;
    mem[4220] = 'd1020;
    mem[4221] = 'd0;
    mem[4222] = 'd1020;
    mem[4223] = 'd0;
    mem[4224] = 'd0;
    mem[4225] = 'd0;
    mem[4226] = 'd1020;
    mem[4227] = 'd0;
    mem[4228] = 'd1020;
    mem[4229] = 'd0;
    mem[4230] = 'd0;
    mem[4231] = 'd0;
    mem[4232] = 'd840;
    mem[4233] = 'd0;
    mem[4234] = 'd924;
    mem[4235] = 'd0;
    mem[4236] = 'd0;
    mem[4237] = 'd0;
    mem[4238] = 'd32;
    mem[4239] = 'd0;
    mem[4240] = 'd608;
    mem[4241] = 'd0;
    mem[4242] = 'd0;
    mem[4243] = 'd0;
    mem[4244] = 'd76;
    mem[4245] = 'd0;
    mem[4246] = 'd736;
    mem[4247] = 'd0;
    mem[4248] = 'd0;
    mem[4249] = 'd0;
    mem[4250] = 'd436;
    mem[4251] = 'd0;
    mem[4252] = 'd896;
    mem[4253] = 'd0;
    mem[4254] = 'd0;
    mem[4255] = 'd0;
    mem[4256] = 'd496;
    mem[4257] = 'd0;
    mem[4258] = 'd936;
    mem[4259] = 'd0;
    mem[4260] = 'd0;
    mem[4261] = 'd0;
    mem[4262] = 'd508;
    mem[4263] = 'd0;
    mem[4264] = 'd956;
    mem[4265] = 'd0;
    mem[4266] = 'd0;
    mem[4267] = 'd0;
    mem[4268] = 'd516;
    mem[4269] = 'd0;
    mem[4270] = 'd976;
    mem[4271] = 'd0;
    mem[4272] = 'd0;
    mem[4273] = 'd0;
    mem[4274] = 'd528;
    mem[4275] = 'd0;
    mem[4276] = 'd992;
    mem[4277] = 'd0;
    mem[4278] = 'd0;
    mem[4279] = 'd0;
    mem[4280] = 'd536;
    mem[4281] = 'd0;
    mem[4282] = 'd992;
    mem[4283] = 'd0;
    mem[4284] = 'd0;
    mem[4285] = 'd0;
    mem[4286] = 'd544;
    mem[4287] = 'd0;
    mem[4288] = 'd996;
    mem[4289] = 'd0;
    mem[4290] = 'd0;
    mem[4291] = 'd0;
    mem[4292] = 'd556;
    mem[4293] = 'd0;
    mem[4294] = 'd996;
    mem[4295] = 'd0;
    mem[4296] = 'd0;
    mem[4297] = 'd0;
    mem[4298] = 'd568;
    mem[4299] = 'd0;
    mem[4300] = 'd996;
    mem[4301] = 'd0;
    mem[4302] = 'd0;
    mem[4303] = 'd0;
    mem[4304] = 'd576;
    mem[4305] = 'd0;
    mem[4306] = 'd996;
    mem[4307] = 'd0;
    mem[4308] = 'd0;
    mem[4309] = 'd0;
    mem[4310] = 'd584;
    mem[4311] = 'd0;
    mem[4312] = 'd996;
    mem[4313] = 'd0;
    mem[4314] = 'd0;
    mem[4315] = 'd0;
    mem[4316] = 'd592;
    mem[4317] = 'd0;
    mem[4318] = 'd996;
    mem[4319] = 'd0;
    mem[4320] = 'd0;
    mem[4321] = 'd0;
    mem[4322] = 'd596;
    mem[4323] = 'd0;
    mem[4324] = 'd996;
    mem[4325] = 'd0;
    mem[4326] = 'd0;
    mem[4327] = 'd0;
    mem[4328] = 'd596;
    mem[4329] = 'd0;
    mem[4330] = 'd996;
    mem[4331] = 'd0;
    mem[4332] = 'd0;
    mem[4333] = 'd0;
    mem[4334] = 'd592;
    mem[4335] = 'd0;
    mem[4336] = 'd996;
    mem[4337] = 'd0;
    mem[4338] = 'd0;
    mem[4339] = 'd0;
    mem[4340] = 'd584;
    mem[4341] = 'd0;
    mem[4342] = 'd996;
    mem[4343] = 'd0;
    mem[4344] = 'd0;
    mem[4345] = 'd0;
    mem[4346] = 'd576;
    mem[4347] = 'd0;
    mem[4348] = 'd996;
    mem[4349] = 'd0;
    mem[4350] = 'd0;
    mem[4351] = 'd0;
    mem[4352] = 'd564;
    mem[4353] = 'd0;
    mem[4354] = 'd996;
    mem[4355] = 'd0;
    mem[4356] = 'd0;
    mem[4357] = 'd0;
    mem[4358] = 'd556;
    mem[4359] = 'd0;
    mem[4360] = 'd996;
    mem[4361] = 'd0;
    mem[4362] = 'd0;
    mem[4363] = 'd0;
    mem[4364] = 'd544;
    mem[4365] = 'd0;
    mem[4366] = 'd996;
    mem[4367] = 'd0;
    mem[4368] = 'd0;
    mem[4369] = 'd0;
    mem[4370] = 'd532;
    mem[4371] = 'd0;
    mem[4372] = 'd992;
    mem[4373] = 'd0;
    mem[4374] = 'd0;
    mem[4375] = 'd0;
    mem[4376] = 'd524;
    mem[4377] = 'd0;
    mem[4378] = 'd992;
    mem[4379] = 'd0;
    mem[4380] = 'd0;
    mem[4381] = 'd0;
    mem[4382] = 'd516;
    mem[4383] = 'd0;
    mem[4384] = 'd976;
    mem[4385] = 'd0;
    mem[4386] = 'd0;
    mem[4387] = 'd0;
    mem[4388] = 'd508;
    mem[4389] = 'd0;
    mem[4390] = 'd956;
    mem[4391] = 'd0;
    mem[4392] = 'd0;
    mem[4393] = 'd0;
    mem[4394] = 'd496;
    mem[4395] = 'd0;
    mem[4396] = 'd936;
    mem[4397] = 'd0;
    mem[4398] = 'd0;
    mem[4399] = 'd0;
    mem[4400] = 'd460;
    mem[4401] = 'd0;
    mem[4402] = 'd900;
    mem[4403] = 'd0;
    mem[4404] = 'd0;
    mem[4405] = 'd0;
    mem[4406] = 'd116;
    mem[4407] = 'd0;
    mem[4408] = 'd748;
    mem[4409] = 'd0;
    mem[4410] = 'd0;
    mem[4411] = 'd0;
    mem[4412] = 'd28;
    mem[4413] = 'd0;
    mem[4414] = 'd604;
    mem[4415] = 'd0;
    mem[4416] = 'd0;
    mem[4417] = 'd0;
    mem[4418] = 'd828;
    mem[4419] = 'd0;
    mem[4420] = 'd912;
    mem[4421] = 'd0;
    mem[4422] = 'd0;
    mem[4423] = 'd0;
    mem[4424] = 'd1020;
    mem[4425] = 'd0;
    mem[4426] = 'd1020;
    mem[4427] = 'd0;
    mem[4428] = 'd0;
    mem[4429] = 'd0;
    mem[4430] = 'd1020;
    mem[4431] = 'd0;
    mem[4432] = 'd1020;
    mem[4433] = 'd0;
    mem[4434] = 'd0;
    mem[4435] = 'd0;
    mem[4436] = 'd1020;
    mem[4437] = 'd0;
    mem[4438] = 'd1020;
    mem[4439] = 'd0;
    mem[4440] = 'd0;
    mem[4441] = 'd0;
    mem[4442] = 'd1020;
    mem[4443] = 'd0;
    mem[4444] = 'd1020;
    mem[4445] = 'd0;
    mem[4446] = 'd0;
    mem[4447] = 'd1020;
    mem[4448] = 'd0;
    mem[4449] = 'd1020;
    mem[4450] = 'd0;
    mem[4451] = 'd0;
    mem[4452] = 'd0;
    mem[4453] = 'd1020;
    mem[4454] = 'd0;
    mem[4455] = 'd1020;
    mem[4456] = 'd0;
    mem[4457] = 'd0;
    mem[4458] = 'd0;
    mem[4459] = 'd1020;
    mem[4460] = 'd0;
    mem[4461] = 'd1020;
    mem[4462] = 'd0;
    mem[4463] = 'd0;
    mem[4464] = 'd0;
    mem[4465] = 'd924;
    mem[4466] = 'd0;
    mem[4467] = 'd996;
    mem[4468] = 'd0;
    mem[4469] = 'd0;
    mem[4470] = 'd0;
    mem[4471] = 'd608;
    mem[4472] = 'd0;
    mem[4473] = 'd1008;
    mem[4474] = 'd0;
    mem[4475] = 'd0;
    mem[4476] = 'd0;
    mem[4477] = 'd736;
    mem[4478] = 'd0;
    mem[4479] = 'd1020;
    mem[4480] = 'd0;
    mem[4481] = 'd0;
    mem[4482] = 'd0;
    mem[4483] = 'd896;
    mem[4484] = 'd0;
    mem[4485] = 'd1020;
    mem[4486] = 'd0;
    mem[4487] = 'd0;
    mem[4488] = 'd0;
    mem[4489] = 'd936;
    mem[4490] = 'd0;
    mem[4491] = 'd1020;
    mem[4492] = 'd0;
    mem[4493] = 'd0;
    mem[4494] = 'd0;
    mem[4495] = 'd956;
    mem[4496] = 'd0;
    mem[4497] = 'd1020;
    mem[4498] = 'd0;
    mem[4499] = 'd0;
    mem[4500] = 'd0;
    mem[4501] = 'd976;
    mem[4502] = 'd0;
    mem[4503] = 'd1020;
    mem[4504] = 'd0;
    mem[4505] = 'd0;
    mem[4506] = 'd0;
    mem[4507] = 'd992;
    mem[4508] = 'd0;
    mem[4509] = 'd1020;
    mem[4510] = 'd0;
    mem[4511] = 'd0;
    mem[4512] = 'd0;
    mem[4513] = 'd992;
    mem[4514] = 'd0;
    mem[4515] = 'd1020;
    mem[4516] = 'd0;
    mem[4517] = 'd0;
    mem[4518] = 'd0;
    mem[4519] = 'd996;
    mem[4520] = 'd0;
    mem[4521] = 'd1020;
    mem[4522] = 'd0;
    mem[4523] = 'd0;
    mem[4524] = 'd0;
    mem[4525] = 'd996;
    mem[4526] = 'd0;
    mem[4527] = 'd1020;
    mem[4528] = 'd0;
    mem[4529] = 'd0;
    mem[4530] = 'd0;
    mem[4531] = 'd996;
    mem[4532] = 'd0;
    mem[4533] = 'd1020;
    mem[4534] = 'd0;
    mem[4535] = 'd0;
    mem[4536] = 'd0;
    mem[4537] = 'd996;
    mem[4538] = 'd0;
    mem[4539] = 'd1020;
    mem[4540] = 'd0;
    mem[4541] = 'd0;
    mem[4542] = 'd0;
    mem[4543] = 'd996;
    mem[4544] = 'd0;
    mem[4545] = 'd1020;
    mem[4546] = 'd0;
    mem[4547] = 'd0;
    mem[4548] = 'd0;
    mem[4549] = 'd996;
    mem[4550] = 'd0;
    mem[4551] = 'd1020;
    mem[4552] = 'd0;
    mem[4553] = 'd0;
    mem[4554] = 'd0;
    mem[4555] = 'd996;
    mem[4556] = 'd0;
    mem[4557] = 'd1020;
    mem[4558] = 'd0;
    mem[4559] = 'd0;
    mem[4560] = 'd0;
    mem[4561] = 'd996;
    mem[4562] = 'd0;
    mem[4563] = 'd1020;
    mem[4564] = 'd0;
    mem[4565] = 'd0;
    mem[4566] = 'd0;
    mem[4567] = 'd996;
    mem[4568] = 'd0;
    mem[4569] = 'd1020;
    mem[4570] = 'd0;
    mem[4571] = 'd0;
    mem[4572] = 'd0;
    mem[4573] = 'd996;
    mem[4574] = 'd0;
    mem[4575] = 'd1020;
    mem[4576] = 'd0;
    mem[4577] = 'd0;
    mem[4578] = 'd0;
    mem[4579] = 'd996;
    mem[4580] = 'd0;
    mem[4581] = 'd1020;
    mem[4582] = 'd0;
    mem[4583] = 'd0;
    mem[4584] = 'd0;
    mem[4585] = 'd996;
    mem[4586] = 'd0;
    mem[4587] = 'd1020;
    mem[4588] = 'd0;
    mem[4589] = 'd0;
    mem[4590] = 'd0;
    mem[4591] = 'd996;
    mem[4592] = 'd0;
    mem[4593] = 'd1020;
    mem[4594] = 'd0;
    mem[4595] = 'd0;
    mem[4596] = 'd0;
    mem[4597] = 'd996;
    mem[4598] = 'd0;
    mem[4599] = 'd1020;
    mem[4600] = 'd0;
    mem[4601] = 'd0;
    mem[4602] = 'd0;
    mem[4603] = 'd992;
    mem[4604] = 'd0;
    mem[4605] = 'd1020;
    mem[4606] = 'd0;
    mem[4607] = 'd0;
    mem[4608] = 'd0;
    mem[4609] = 'd992;
    mem[4610] = 'd0;
    mem[4611] = 'd1020;
    mem[4612] = 'd0;
    mem[4613] = 'd0;
    mem[4614] = 'd0;
    mem[4615] = 'd976;
    mem[4616] = 'd0;
    mem[4617] = 'd1020;
    mem[4618] = 'd0;
    mem[4619] = 'd0;
    mem[4620] = 'd0;
    mem[4621] = 'd956;
    mem[4622] = 'd0;
    mem[4623] = 'd1020;
    mem[4624] = 'd0;
    mem[4625] = 'd0;
    mem[4626] = 'd0;
    mem[4627] = 'd936;
    mem[4628] = 'd0;
    mem[4629] = 'd1020;
    mem[4630] = 'd0;
    mem[4631] = 'd0;
    mem[4632] = 'd0;
    mem[4633] = 'd900;
    mem[4634] = 'd0;
    mem[4635] = 'd1020;
    mem[4636] = 'd0;
    mem[4637] = 'd0;
    mem[4638] = 'd0;
    mem[4639] = 'd748;
    mem[4640] = 'd0;
    mem[4641] = 'd1020;
    mem[4642] = 'd0;
    mem[4643] = 'd0;
    mem[4644] = 'd0;
    mem[4645] = 'd604;
    mem[4646] = 'd0;
    mem[4647] = 'd1012;
    mem[4648] = 'd0;
    mem[4649] = 'd0;
    mem[4650] = 'd0;
    mem[4651] = 'd912;
    mem[4652] = 'd0;
    mem[4653] = 'd988;
    mem[4654] = 'd0;
    mem[4655] = 'd0;
    mem[4656] = 'd0;
    mem[4657] = 'd1020;
    mem[4658] = 'd0;
    mem[4659] = 'd1020;
    mem[4660] = 'd0;
    mem[4661] = 'd0;
    mem[4662] = 'd0;
    mem[4663] = 'd1020;
    mem[4664] = 'd0;
    mem[4665] = 'd1020;
    mem[4666] = 'd0;
    mem[4667] = 'd0;
    mem[4668] = 'd0;
    mem[4669] = 'd1020;
    mem[4670] = 'd0;
    mem[4671] = 'd1020;
    mem[4672] = 'd0;
    mem[4673] = 'd0;
    mem[4674] = 'd0;
    mem[4675] = 'd1020;
    mem[4676] = 'd0;
    mem[4677] = 'd1020;
    mem[4678] = 'd0;
    mem[4679] = 'd0;
    mem[4680] = 'd0;
    mem[4681] = 'd0;
    mem[4682] = 'd1020;
    mem[4683] = 'd0;
    mem[4684] = 'd1020;
    mem[4685] = 'd0;
    mem[4686] = 'd0;
    mem[4687] = 'd0;
    mem[4688] = 'd1020;
    mem[4689] = 'd0;
    mem[4690] = 'd1020;
    mem[4691] = 'd0;
    mem[4692] = 'd0;
    mem[4693] = 'd0;
    mem[4694] = 'd1012;
    mem[4695] = 'd0;
    mem[4696] = 'd1016;
    mem[4697] = 'd0;
    mem[4698] = 'd0;
    mem[4699] = 'd0;
    mem[4700] = 'd304;
    mem[4701] = 'd0;
    mem[4702] = 'd668;
    mem[4703] = 'd0;
    mem[4704] = 'd0;
    mem[4705] = 'd0;
    mem[4706] = 'd32;
    mem[4707] = 'd0;
    mem[4708] = 'd668;
    mem[4709] = 'd0;
    mem[4710] = 'd0;
    mem[4711] = 'd0;
    mem[4712] = 'd284;
    mem[4713] = 'd0;
    mem[4714] = 'd824;
    mem[4715] = 'd0;
    mem[4716] = 'd0;
    mem[4717] = 'd0;
    mem[4718] = 'd428;
    mem[4719] = 'd0;
    mem[4720] = 'd900;
    mem[4721] = 'd0;
    mem[4722] = 'd0;
    mem[4723] = 'd0;
    mem[4724] = 'd440;
    mem[4725] = 'd0;
    mem[4726] = 'd924;
    mem[4727] = 'd0;
    mem[4728] = 'd0;
    mem[4729] = 'd0;
    mem[4730] = 'd452;
    mem[4731] = 'd0;
    mem[4732] = 'd948;
    mem[4733] = 'd0;
    mem[4734] = 'd0;
    mem[4735] = 'd0;
    mem[4736] = 'd456;
    mem[4737] = 'd0;
    mem[4738] = 'd964;
    mem[4739] = 'd0;
    mem[4740] = 'd0;
    mem[4741] = 'd0;
    mem[4742] = 'd464;
    mem[4743] = 'd0;
    mem[4744] = 'd976;
    mem[4745] = 'd0;
    mem[4746] = 'd0;
    mem[4747] = 'd0;
    mem[4748] = 'd476;
    mem[4749] = 'd0;
    mem[4750] = 'd988;
    mem[4751] = 'd0;
    mem[4752] = 'd0;
    mem[4753] = 'd0;
    mem[4754] = 'd484;
    mem[4755] = 'd0;
    mem[4756] = 'd988;
    mem[4757] = 'd0;
    mem[4758] = 'd0;
    mem[4759] = 'd0;
    mem[4760] = 'd492;
    mem[4761] = 'd0;
    mem[4762] = 'd988;
    mem[4763] = 'd0;
    mem[4764] = 'd0;
    mem[4765] = 'd0;
    mem[4766] = 'd504;
    mem[4767] = 'd0;
    mem[4768] = 'd992;
    mem[4769] = 'd0;
    mem[4770] = 'd0;
    mem[4771] = 'd0;
    mem[4772] = 'd512;
    mem[4773] = 'd0;
    mem[4774] = 'd992;
    mem[4775] = 'd0;
    mem[4776] = 'd0;
    mem[4777] = 'd0;
    mem[4778] = 'd520;
    mem[4779] = 'd0;
    mem[4780] = 'd992;
    mem[4781] = 'd0;
    mem[4782] = 'd0;
    mem[4783] = 'd0;
    mem[4784] = 'd524;
    mem[4785] = 'd0;
    mem[4786] = 'd992;
    mem[4787] = 'd0;
    mem[4788] = 'd0;
    mem[4789] = 'd0;
    mem[4790] = 'd528;
    mem[4791] = 'd0;
    mem[4792] = 'd992;
    mem[4793] = 'd0;
    mem[4794] = 'd0;
    mem[4795] = 'd0;
    mem[4796] = 'd528;
    mem[4797] = 'd0;
    mem[4798] = 'd992;
    mem[4799] = 'd0;
    mem[4800] = 'd0;
    mem[4801] = 'd0;
    mem[4802] = 'd524;
    mem[4803] = 'd0;
    mem[4804] = 'd992;
    mem[4805] = 'd0;
    mem[4806] = 'd0;
    mem[4807] = 'd0;
    mem[4808] = 'd520;
    mem[4809] = 'd0;
    mem[4810] = 'd992;
    mem[4811] = 'd0;
    mem[4812] = 'd0;
    mem[4813] = 'd0;
    mem[4814] = 'd508;
    mem[4815] = 'd0;
    mem[4816] = 'd992;
    mem[4817] = 'd0;
    mem[4818] = 'd0;
    mem[4819] = 'd0;
    mem[4820] = 'd504;
    mem[4821] = 'd0;
    mem[4822] = 'd992;
    mem[4823] = 'd0;
    mem[4824] = 'd0;
    mem[4825] = 'd0;
    mem[4826] = 'd492;
    mem[4827] = 'd0;
    mem[4828] = 'd988;
    mem[4829] = 'd0;
    mem[4830] = 'd0;
    mem[4831] = 'd0;
    mem[4832] = 'd484;
    mem[4833] = 'd0;
    mem[4834] = 'd988;
    mem[4835] = 'd0;
    mem[4836] = 'd0;
    mem[4837] = 'd0;
    mem[4838] = 'd476;
    mem[4839] = 'd0;
    mem[4840] = 'd988;
    mem[4841] = 'd0;
    mem[4842] = 'd0;
    mem[4843] = 'd0;
    mem[4844] = 'd464;
    mem[4845] = 'd0;
    mem[4846] = 'd976;
    mem[4847] = 'd0;
    mem[4848] = 'd0;
    mem[4849] = 'd0;
    mem[4850] = 'd460;
    mem[4851] = 'd0;
    mem[4852] = 'd964;
    mem[4853] = 'd0;
    mem[4854] = 'd0;
    mem[4855] = 'd0;
    mem[4856] = 'd448;
    mem[4857] = 'd0;
    mem[4858] = 'd948;
    mem[4859] = 'd0;
    mem[4860] = 'd0;
    mem[4861] = 'd0;
    mem[4862] = 'd440;
    mem[4863] = 'd0;
    mem[4864] = 'd928;
    mem[4865] = 'd0;
    mem[4866] = 'd0;
    mem[4867] = 'd0;
    mem[4868] = 'd428;
    mem[4869] = 'd0;
    mem[4870] = 'd900;
    mem[4871] = 'd0;
    mem[4872] = 'd0;
    mem[4873] = 'd0;
    mem[4874] = 'd336;
    mem[4875] = 'd0;
    mem[4876] = 'd844;
    mem[4877] = 'd0;
    mem[4878] = 'd0;
    mem[4879] = 'd0;
    mem[4880] = 'd40;
    mem[4881] = 'd0;
    mem[4882] = 'd672;
    mem[4883] = 'd0;
    mem[4884] = 'd0;
    mem[4885] = 'd0;
    mem[4886] = 'd256;
    mem[4887] = 'd0;
    mem[4888] = 'd644;
    mem[4889] = 'd0;
    mem[4890] = 'd0;
    mem[4891] = 'd0;
    mem[4892] = 'd1020;
    mem[4893] = 'd0;
    mem[4894] = 'd1020;
    mem[4895] = 'd0;
    mem[4896] = 'd0;
    mem[4897] = 'd0;
    mem[4898] = 'd1020;
    mem[4899] = 'd0;
    mem[4900] = 'd1020;
    mem[4901] = 'd0;
    mem[4902] = 'd0;
    mem[4903] = 'd0;
    mem[4904] = 'd1020;
    mem[4905] = 'd0;
    mem[4906] = 'd1020;
    mem[4907] = 'd0;
    mem[4908] = 'd0;
    mem[4909] = 'd0;
    mem[4910] = 'd1020;
    mem[4911] = 'd0;
    mem[4912] = 'd1020;
    mem[4913] = 'd0;
    mem[4914] = 'd0;
    mem[4915] = 'd1020;
    mem[4916] = 'd0;
    mem[4917] = 'd1020;
    mem[4918] = 'd0;
    mem[4919] = 'd0;
    mem[4920] = 'd0;
    mem[4921] = 'd1020;
    mem[4922] = 'd0;
    mem[4923] = 'd1020;
    mem[4924] = 'd0;
    mem[4925] = 'd0;
    mem[4926] = 'd0;
    mem[4927] = 'd1016;
    mem[4928] = 'd0;
    mem[4929] = 'd1016;
    mem[4930] = 'd0;
    mem[4931] = 'd0;
    mem[4932] = 'd0;
    mem[4933] = 'd668;
    mem[4934] = 'd0;
    mem[4935] = 'd972;
    mem[4936] = 'd0;
    mem[4937] = 'd0;
    mem[4938] = 'd0;
    mem[4939] = 'd668;
    mem[4940] = 'd0;
    mem[4941] = 'd1020;
    mem[4942] = 'd0;
    mem[4943] = 'd0;
    mem[4944] = 'd0;
    mem[4945] = 'd824;
    mem[4946] = 'd0;
    mem[4947] = 'd1020;
    mem[4948] = 'd0;
    mem[4949] = 'd0;
    mem[4950] = 'd0;
    mem[4951] = 'd900;
    mem[4952] = 'd0;
    mem[4953] = 'd1020;
    mem[4954] = 'd0;
    mem[4955] = 'd0;
    mem[4956] = 'd0;
    mem[4957] = 'd924;
    mem[4958] = 'd0;
    mem[4959] = 'd1020;
    mem[4960] = 'd0;
    mem[4961] = 'd0;
    mem[4962] = 'd0;
    mem[4963] = 'd948;
    mem[4964] = 'd0;
    mem[4965] = 'd1020;
    mem[4966] = 'd0;
    mem[4967] = 'd0;
    mem[4968] = 'd0;
    mem[4969] = 'd964;
    mem[4970] = 'd0;
    mem[4971] = 'd1020;
    mem[4972] = 'd0;
    mem[4973] = 'd0;
    mem[4974] = 'd0;
    mem[4975] = 'd976;
    mem[4976] = 'd0;
    mem[4977] = 'd1020;
    mem[4978] = 'd0;
    mem[4979] = 'd0;
    mem[4980] = 'd0;
    mem[4981] = 'd988;
    mem[4982] = 'd0;
    mem[4983] = 'd1020;
    mem[4984] = 'd0;
    mem[4985] = 'd0;
    mem[4986] = 'd0;
    mem[4987] = 'd988;
    mem[4988] = 'd0;
    mem[4989] = 'd1020;
    mem[4990] = 'd0;
    mem[4991] = 'd0;
    mem[4992] = 'd0;
    mem[4993] = 'd988;
    mem[4994] = 'd0;
    mem[4995] = 'd1020;
    mem[4996] = 'd0;
    mem[4997] = 'd0;
    mem[4998] = 'd0;
    mem[4999] = 'd992;
    mem[5000] = 'd0;
    mem[5001] = 'd1020;
    mem[5002] = 'd0;
    mem[5003] = 'd0;
    mem[5004] = 'd0;
    mem[5005] = 'd992;
    mem[5006] = 'd0;
    mem[5007] = 'd1020;
    mem[5008] = 'd0;
    mem[5009] = 'd0;
    mem[5010] = 'd0;
    mem[5011] = 'd992;
    mem[5012] = 'd0;
    mem[5013] = 'd1020;
    mem[5014] = 'd0;
    mem[5015] = 'd0;
    mem[5016] = 'd0;
    mem[5017] = 'd992;
    mem[5018] = 'd0;
    mem[5019] = 'd1020;
    mem[5020] = 'd0;
    mem[5021] = 'd0;
    mem[5022] = 'd0;
    mem[5023] = 'd992;
    mem[5024] = 'd0;
    mem[5025] = 'd1020;
    mem[5026] = 'd0;
    mem[5027] = 'd0;
    mem[5028] = 'd0;
    mem[5029] = 'd992;
    mem[5030] = 'd0;
    mem[5031] = 'd1020;
    mem[5032] = 'd0;
    mem[5033] = 'd0;
    mem[5034] = 'd0;
    mem[5035] = 'd992;
    mem[5036] = 'd0;
    mem[5037] = 'd1020;
    mem[5038] = 'd0;
    mem[5039] = 'd0;
    mem[5040] = 'd0;
    mem[5041] = 'd992;
    mem[5042] = 'd0;
    mem[5043] = 'd1020;
    mem[5044] = 'd0;
    mem[5045] = 'd0;
    mem[5046] = 'd0;
    mem[5047] = 'd992;
    mem[5048] = 'd0;
    mem[5049] = 'd1020;
    mem[5050] = 'd0;
    mem[5051] = 'd0;
    mem[5052] = 'd0;
    mem[5053] = 'd992;
    mem[5054] = 'd0;
    mem[5055] = 'd1020;
    mem[5056] = 'd0;
    mem[5057] = 'd0;
    mem[5058] = 'd0;
    mem[5059] = 'd988;
    mem[5060] = 'd0;
    mem[5061] = 'd1020;
    mem[5062] = 'd0;
    mem[5063] = 'd0;
    mem[5064] = 'd0;
    mem[5065] = 'd988;
    mem[5066] = 'd0;
    mem[5067] = 'd1020;
    mem[5068] = 'd0;
    mem[5069] = 'd0;
    mem[5070] = 'd0;
    mem[5071] = 'd988;
    mem[5072] = 'd0;
    mem[5073] = 'd1020;
    mem[5074] = 'd0;
    mem[5075] = 'd0;
    mem[5076] = 'd0;
    mem[5077] = 'd976;
    mem[5078] = 'd0;
    mem[5079] = 'd1020;
    mem[5080] = 'd0;
    mem[5081] = 'd0;
    mem[5082] = 'd0;
    mem[5083] = 'd964;
    mem[5084] = 'd0;
    mem[5085] = 'd1020;
    mem[5086] = 'd0;
    mem[5087] = 'd0;
    mem[5088] = 'd0;
    mem[5089] = 'd948;
    mem[5090] = 'd0;
    mem[5091] = 'd1020;
    mem[5092] = 'd0;
    mem[5093] = 'd0;
    mem[5094] = 'd0;
    mem[5095] = 'd928;
    mem[5096] = 'd0;
    mem[5097] = 'd1020;
    mem[5098] = 'd0;
    mem[5099] = 'd0;
    mem[5100] = 'd0;
    mem[5101] = 'd900;
    mem[5102] = 'd0;
    mem[5103] = 'd1020;
    mem[5104] = 'd0;
    mem[5105] = 'd0;
    mem[5106] = 'd0;
    mem[5107] = 'd844;
    mem[5108] = 'd0;
    mem[5109] = 'd1020;
    mem[5110] = 'd0;
    mem[5111] = 'd0;
    mem[5112] = 'd0;
    mem[5113] = 'd672;
    mem[5114] = 'd0;
    mem[5115] = 'd1020;
    mem[5116] = 'd0;
    mem[5117] = 'd0;
    mem[5118] = 'd0;
    mem[5119] = 'd644;
    mem[5120] = 'd0;
    mem[5121] = 'd972;
    mem[5122] = 'd0;
    mem[5123] = 'd0;
    mem[5124] = 'd0;
    mem[5125] = 'd1020;
    mem[5126] = 'd0;
    mem[5127] = 'd1020;
    mem[5128] = 'd0;
    mem[5129] = 'd0;
    mem[5130] = 'd0;
    mem[5131] = 'd1020;
    mem[5132] = 'd0;
    mem[5133] = 'd1020;
    mem[5134] = 'd0;
    mem[5135] = 'd0;
    mem[5136] = 'd0;
    mem[5137] = 'd1020;
    mem[5138] = 'd0;
    mem[5139] = 'd1020;
    mem[5140] = 'd0;
    mem[5141] = 'd0;
    mem[5142] = 'd0;
    mem[5143] = 'd1020;
    mem[5144] = 'd0;
    mem[5145] = 'd1020;
    mem[5146] = 'd0;
    mem[5147] = 'd0;
    mem[5148] = 'd0;
    mem[5149] = 'd0;
    mem[5150] = 'd1020;
    mem[5151] = 'd0;
    mem[5152] = 'd1020;
    mem[5153] = 'd0;
    mem[5154] = 'd0;
    mem[5155] = 'd0;
    mem[5156] = 'd1020;
    mem[5157] = 'd0;
    mem[5158] = 'd1020;
    mem[5159] = 'd0;
    mem[5160] = 'd0;
    mem[5161] = 'd0;
    mem[5162] = 'd788;
    mem[5163] = 'd0;
    mem[5164] = 'd892;
    mem[5165] = 'd0;
    mem[5166] = 'd0;
    mem[5167] = 'd0;
    mem[5168] = 'd24;
    mem[5169] = 'd0;
    mem[5170] = 'd584;
    mem[5171] = 'd0;
    mem[5172] = 'd0;
    mem[5173] = 'd0;
    mem[5174] = 'd108;
    mem[5175] = 'd0;
    mem[5176] = 'd700;
    mem[5177] = 'd0;
    mem[5178] = 'd0;
    mem[5179] = 'd0;
    mem[5180] = 'd344;
    mem[5181] = 'd0;
    mem[5182] = 'd804;
    mem[5183] = 'd0;
    mem[5184] = 'd0;
    mem[5185] = 'd0;
    mem[5186] = 'd356;
    mem[5187] = 'd0;
    mem[5188] = 'd824;
    mem[5189] = 'd0;
    mem[5190] = 'd0;
    mem[5191] = 'd0;
    mem[5192] = 'd364;
    mem[5193] = 'd0;
    mem[5194] = 'd840;
    mem[5195] = 'd0;
    mem[5196] = 'd0;
    mem[5197] = 'd0;
    mem[5198] = 'd372;
    mem[5199] = 'd0;
    mem[5200] = 'd860;
    mem[5201] = 'd0;
    mem[5202] = 'd0;
    mem[5203] = 'd0;
    mem[5204] = 'd388;
    mem[5205] = 'd0;
    mem[5206] = 'd888;
    mem[5207] = 'd0;
    mem[5208] = 'd0;
    mem[5209] = 'd0;
    mem[5210] = 'd396;
    mem[5211] = 'd0;
    mem[5212] = 'd912;
    mem[5213] = 'd0;
    mem[5214] = 'd0;
    mem[5215] = 'd0;
    mem[5216] = 'd408;
    mem[5217] = 'd0;
    mem[5218] = 'd952;
    mem[5219] = 'd0;
    mem[5220] = 'd0;
    mem[5221] = 'd0;
    mem[5222] = 'd424;
    mem[5223] = 'd0;
    mem[5224] = 'd988;
    mem[5225] = 'd0;
    mem[5226] = 'd0;
    mem[5227] = 'd0;
    mem[5228] = 'd436;
    mem[5229] = 'd0;
    mem[5230] = 'd992;
    mem[5231] = 'd0;
    mem[5232] = 'd0;
    mem[5233] = 'd0;
    mem[5234] = 'd436;
    mem[5235] = 'd0;
    mem[5236] = 'd988;
    mem[5237] = 'd0;
    mem[5238] = 'd0;
    mem[5239] = 'd0;
    mem[5240] = 'd448;
    mem[5241] = 'd0;
    mem[5242] = 'd988;
    mem[5243] = 'd0;
    mem[5244] = 'd0;
    mem[5245] = 'd0;
    mem[5246] = 'd456;
    mem[5247] = 'd0;
    mem[5248] = 'd988;
    mem[5249] = 'd0;
    mem[5250] = 'd0;
    mem[5251] = 'd0;
    mem[5252] = 'd456;
    mem[5253] = 'd0;
    mem[5254] = 'd988;
    mem[5255] = 'd0;
    mem[5256] = 'd0;
    mem[5257] = 'd0;
    mem[5258] = 'd460;
    mem[5259] = 'd0;
    mem[5260] = 'd988;
    mem[5261] = 'd0;
    mem[5262] = 'd0;
    mem[5263] = 'd0;
    mem[5264] = 'd460;
    mem[5265] = 'd0;
    mem[5266] = 'd988;
    mem[5267] = 'd0;
    mem[5268] = 'd0;
    mem[5269] = 'd0;
    mem[5270] = 'd460;
    mem[5271] = 'd0;
    mem[5272] = 'd988;
    mem[5273] = 'd0;
    mem[5274] = 'd0;
    mem[5275] = 'd0;
    mem[5276] = 'd456;
    mem[5277] = 'd0;
    mem[5278] = 'd988;
    mem[5279] = 'd0;
    mem[5280] = 'd0;
    mem[5281] = 'd0;
    mem[5282] = 'd444;
    mem[5283] = 'd0;
    mem[5284] = 'd988;
    mem[5285] = 'd0;
    mem[5286] = 'd0;
    mem[5287] = 'd0;
    mem[5288] = 'd436;
    mem[5289] = 'd0;
    mem[5290] = 'd992;
    mem[5291] = 'd0;
    mem[5292] = 'd0;
    mem[5293] = 'd0;
    mem[5294] = 'd432;
    mem[5295] = 'd0;
    mem[5296] = 'd992;
    mem[5297] = 'd0;
    mem[5298] = 'd0;
    mem[5299] = 'd0;
    mem[5300] = 'd424;
    mem[5301] = 'd0;
    mem[5302] = 'd980;
    mem[5303] = 'd0;
    mem[5304] = 'd0;
    mem[5305] = 'd0;
    mem[5306] = 'd404;
    mem[5307] = 'd0;
    mem[5308] = 'd944;
    mem[5309] = 'd0;
    mem[5310] = 'd0;
    mem[5311] = 'd0;
    mem[5312] = 'd392;
    mem[5313] = 'd0;
    mem[5314] = 'd908;
    mem[5315] = 'd0;
    mem[5316] = 'd0;
    mem[5317] = 'd0;
    mem[5318] = 'd380;
    mem[5319] = 'd0;
    mem[5320] = 'd884;
    mem[5321] = 'd0;
    mem[5322] = 'd0;
    mem[5323] = 'd0;
    mem[5324] = 'd376;
    mem[5325] = 'd0;
    mem[5326] = 'd860;
    mem[5327] = 'd0;
    mem[5328] = 'd0;
    mem[5329] = 'd0;
    mem[5330] = 'd368;
    mem[5331] = 'd0;
    mem[5332] = 'd844;
    mem[5333] = 'd0;
    mem[5334] = 'd0;
    mem[5335] = 'd0;
    mem[5336] = 'd356;
    mem[5337] = 'd0;
    mem[5338] = 'd828;
    mem[5339] = 'd0;
    mem[5340] = 'd0;
    mem[5341] = 'd0;
    mem[5342] = 'd348;
    mem[5343] = 'd0;
    mem[5344] = 'd812;
    mem[5345] = 'd0;
    mem[5346] = 'd0;
    mem[5347] = 'd0;
    mem[5348] = 'd148;
    mem[5349] = 'd0;
    mem[5350] = 'd728;
    mem[5351] = 'd0;
    mem[5352] = 'd0;
    mem[5353] = 'd0;
    mem[5354] = 'd16;
    mem[5355] = 'd0;
    mem[5356] = 'd584;
    mem[5357] = 'd0;
    mem[5358] = 'd0;
    mem[5359] = 'd0;
    mem[5360] = 'd760;
    mem[5361] = 'd0;
    mem[5362] = 'd872;
    mem[5363] = 'd0;
    mem[5364] = 'd0;
    mem[5365] = 'd0;
    mem[5366] = 'd1020;
    mem[5367] = 'd0;
    mem[5368] = 'd1020;
    mem[5369] = 'd0;
    mem[5370] = 'd0;
    mem[5371] = 'd0;
    mem[5372] = 'd1020;
    mem[5373] = 'd0;
    mem[5374] = 'd1020;
    mem[5375] = 'd0;
    mem[5376] = 'd0;
    mem[5377] = 'd0;
    mem[5378] = 'd1020;
    mem[5379] = 'd0;
    mem[5380] = 'd1020;
    mem[5381] = 'd0;
    mem[5382] = 'd0;
    mem[5383] = 'd1020;
    mem[5384] = 'd0;
    mem[5385] = 'd1020;
    mem[5386] = 'd0;
    mem[5387] = 'd0;
    mem[5388] = 'd0;
    mem[5389] = 'd1020;
    mem[5390] = 'd0;
    mem[5391] = 'd1020;
    mem[5392] = 'd0;
    mem[5393] = 'd0;
    mem[5394] = 'd0;
    mem[5395] = 'd892;
    mem[5396] = 'd0;
    mem[5397] = 'd984;
    mem[5398] = 'd0;
    mem[5399] = 'd0;
    mem[5400] = 'd0;
    mem[5401] = 'd584;
    mem[5402] = 'd0;
    mem[5403] = 'd1000;
    mem[5404] = 'd0;
    mem[5405] = 'd0;
    mem[5406] = 'd0;
    mem[5407] = 'd700;
    mem[5408] = 'd0;
    mem[5409] = 'd968;
    mem[5410] = 'd0;
    mem[5411] = 'd0;
    mem[5412] = 'd0;
    mem[5413] = 'd804;
    mem[5414] = 'd0;
    mem[5415] = 'd948;
    mem[5416] = 'd0;
    mem[5417] = 'd0;
    mem[5418] = 'd0;
    mem[5419] = 'd824;
    mem[5420] = 'd0;
    mem[5421] = 'd940;
    mem[5422] = 'd0;
    mem[5423] = 'd0;
    mem[5424] = 'd0;
    mem[5425] = 'd840;
    mem[5426] = 'd0;
    mem[5427] = 'd932;
    mem[5428] = 'd0;
    mem[5429] = 'd0;
    mem[5430] = 'd0;
    mem[5431] = 'd860;
    mem[5432] = 'd0;
    mem[5433] = 'd936;
    mem[5434] = 'd0;
    mem[5435] = 'd0;
    mem[5436] = 'd0;
    mem[5437] = 'd888;
    mem[5438] = 'd0;
    mem[5439] = 'd944;
    mem[5440] = 'd0;
    mem[5441] = 'd0;
    mem[5442] = 'd0;
    mem[5443] = 'd912;
    mem[5444] = 'd0;
    mem[5445] = 'd956;
    mem[5446] = 'd0;
    mem[5447] = 'd0;
    mem[5448] = 'd0;
    mem[5449] = 'd952;
    mem[5450] = 'd0;
    mem[5451] = 'd980;
    mem[5452] = 'd0;
    mem[5453] = 'd0;
    mem[5454] = 'd0;
    mem[5455] = 'd988;
    mem[5456] = 'd0;
    mem[5457] = 'd1012;
    mem[5458] = 'd0;
    mem[5459] = 'd0;
    mem[5460] = 'd0;
    mem[5461] = 'd992;
    mem[5462] = 'd0;
    mem[5463] = 'd1020;
    mem[5464] = 'd0;
    mem[5465] = 'd0;
    mem[5466] = 'd0;
    mem[5467] = 'd988;
    mem[5468] = 'd0;
    mem[5469] = 'd1020;
    mem[5470] = 'd0;
    mem[5471] = 'd0;
    mem[5472] = 'd0;
    mem[5473] = 'd988;
    mem[5474] = 'd0;
    mem[5475] = 'd1020;
    mem[5476] = 'd0;
    mem[5477] = 'd0;
    mem[5478] = 'd0;
    mem[5479] = 'd988;
    mem[5480] = 'd0;
    mem[5481] = 'd1020;
    mem[5482] = 'd0;
    mem[5483] = 'd0;
    mem[5484] = 'd0;
    mem[5485] = 'd988;
    mem[5486] = 'd0;
    mem[5487] = 'd1020;
    mem[5488] = 'd0;
    mem[5489] = 'd0;
    mem[5490] = 'd0;
    mem[5491] = 'd988;
    mem[5492] = 'd0;
    mem[5493] = 'd1020;
    mem[5494] = 'd0;
    mem[5495] = 'd0;
    mem[5496] = 'd0;
    mem[5497] = 'd988;
    mem[5498] = 'd0;
    mem[5499] = 'd1020;
    mem[5500] = 'd0;
    mem[5501] = 'd0;
    mem[5502] = 'd0;
    mem[5503] = 'd988;
    mem[5504] = 'd0;
    mem[5505] = 'd1020;
    mem[5506] = 'd0;
    mem[5507] = 'd0;
    mem[5508] = 'd0;
    mem[5509] = 'd988;
    mem[5510] = 'd0;
    mem[5511] = 'd1020;
    mem[5512] = 'd0;
    mem[5513] = 'd0;
    mem[5514] = 'd0;
    mem[5515] = 'd988;
    mem[5516] = 'd0;
    mem[5517] = 'd1020;
    mem[5518] = 'd0;
    mem[5519] = 'd0;
    mem[5520] = 'd0;
    mem[5521] = 'd992;
    mem[5522] = 'd0;
    mem[5523] = 'd1020;
    mem[5524] = 'd0;
    mem[5525] = 'd0;
    mem[5526] = 'd0;
    mem[5527] = 'd992;
    mem[5528] = 'd0;
    mem[5529] = 'd1020;
    mem[5530] = 'd0;
    mem[5531] = 'd0;
    mem[5532] = 'd0;
    mem[5533] = 'd980;
    mem[5534] = 'd0;
    mem[5535] = 'd1008;
    mem[5536] = 'd0;
    mem[5537] = 'd0;
    mem[5538] = 'd0;
    mem[5539] = 'd944;
    mem[5540] = 'd0;
    mem[5541] = 'd976;
    mem[5542] = 'd0;
    mem[5543] = 'd0;
    mem[5544] = 'd0;
    mem[5545] = 'd908;
    mem[5546] = 'd0;
    mem[5547] = 'd956;
    mem[5548] = 'd0;
    mem[5549] = 'd0;
    mem[5550] = 'd0;
    mem[5551] = 'd884;
    mem[5552] = 'd0;
    mem[5553] = 'd940;
    mem[5554] = 'd0;
    mem[5555] = 'd0;
    mem[5556] = 'd0;
    mem[5557] = 'd860;
    mem[5558] = 'd0;
    mem[5559] = 'd932;
    mem[5560] = 'd0;
    mem[5561] = 'd0;
    mem[5562] = 'd0;
    mem[5563] = 'd844;
    mem[5564] = 'd0;
    mem[5565] = 'd936;
    mem[5566] = 'd0;
    mem[5567] = 'd0;
    mem[5568] = 'd0;
    mem[5569] = 'd828;
    mem[5570] = 'd0;
    mem[5571] = 'd940;
    mem[5572] = 'd0;
    mem[5573] = 'd0;
    mem[5574] = 'd0;
    mem[5575] = 'd812;
    mem[5576] = 'd0;
    mem[5577] = 'd952;
    mem[5578] = 'd0;
    mem[5579] = 'd0;
    mem[5580] = 'd0;
    mem[5581] = 'd728;
    mem[5582] = 'd0;
    mem[5583] = 'd988;
    mem[5584] = 'd0;
    mem[5585] = 'd0;
    mem[5586] = 'd0;
    mem[5587] = 'd584;
    mem[5588] = 'd0;
    mem[5589] = 'd1004;
    mem[5590] = 'd0;
    mem[5591] = 'd0;
    mem[5592] = 'd0;
    mem[5593] = 'd872;
    mem[5594] = 'd0;
    mem[5595] = 'd976;
    mem[5596] = 'd0;
    mem[5597] = 'd0;
    mem[5598] = 'd0;
    mem[5599] = 'd1020;
    mem[5600] = 'd0;
    mem[5601] = 'd1020;
    mem[5602] = 'd0;
    mem[5603] = 'd0;
    mem[5604] = 'd0;
    mem[5605] = 'd1020;
    mem[5606] = 'd0;
    mem[5607] = 'd1020;
    mem[5608] = 'd0;
    mem[5609] = 'd0;
    mem[5610] = 'd0;
    mem[5611] = 'd1020;
    mem[5612] = 'd0;
    mem[5613] = 'd1020;
    mem[5614] = 'd0;
    mem[5615] = 'd0;
    mem[5616] = 'd0;
    mem[5617] = 'd0;
    mem[5618] = 'd1020;
    mem[5619] = 'd0;
    mem[5620] = 'd1020;
    mem[5621] = 'd0;
    mem[5622] = 'd0;
    mem[5623] = 'd0;
    mem[5624] = 'd1020;
    mem[5625] = 'd0;
    mem[5626] = 'd1020;
    mem[5627] = 'd0;
    mem[5628] = 'd0;
    mem[5629] = 'd0;
    mem[5630] = 'd352;
    mem[5631] = 'd0;
    mem[5632] = 'd676;
    mem[5633] = 'd0;
    mem[5634] = 'd0;
    mem[5635] = 'd0;
    mem[5636] = 'd52;
    mem[5637] = 'd0;
    mem[5638] = 'd460;
    mem[5639] = 'd0;
    mem[5640] = 'd0;
    mem[5641] = 'd0;
    mem[5642] = 'd132;
    mem[5643] = 'd0;
    mem[5644] = 'd168;
    mem[5645] = 'd0;
    mem[5646] = 'd0;
    mem[5647] = 'd0;
    mem[5648] = 'd152;
    mem[5649] = 'd0;
    mem[5650] = 'd168;
    mem[5651] = 'd0;
    mem[5652] = 'd0;
    mem[5653] = 'd0;
    mem[5654] = 'd152;
    mem[5655] = 'd0;
    mem[5656] = 'd168;
    mem[5657] = 'd0;
    mem[5658] = 'd0;
    mem[5659] = 'd0;
    mem[5660] = 'd148;
    mem[5661] = 'd0;
    mem[5662] = 'd160;
    mem[5663] = 'd0;
    mem[5664] = 'd0;
    mem[5665] = 'd0;
    mem[5666] = 'd140;
    mem[5667] = 'd0;
    mem[5668] = 'd152;
    mem[5669] = 'd0;
    mem[5670] = 'd0;
    mem[5671] = 'd0;
    mem[5672] = 'd144;
    mem[5673] = 'd0;
    mem[5674] = 'd160;
    mem[5675] = 'd0;
    mem[5676] = 'd0;
    mem[5677] = 'd0;
    mem[5678] = 'd152;
    mem[5679] = 'd0;
    mem[5680] = 'd176;
    mem[5681] = 'd0;
    mem[5682] = 'd0;
    mem[5683] = 'd0;
    mem[5684] = 'd172;
    mem[5685] = 'd0;
    mem[5686] = 'd220;
    mem[5687] = 'd0;
    mem[5688] = 'd0;
    mem[5689] = 'd0;
    mem[5690] = 'd204;
    mem[5691] = 'd0;
    mem[5692] = 'd304;
    mem[5693] = 'd0;
    mem[5694] = 'd0;
    mem[5695] = 'd0;
    mem[5696] = 'd248;
    mem[5697] = 'd0;
    mem[5698] = 'd428;
    mem[5699] = 'd0;
    mem[5700] = 'd0;
    mem[5701] = 'd0;
    mem[5702] = 'd308;
    mem[5703] = 'd0;
    mem[5704] = 'd628;
    mem[5705] = 'd0;
    mem[5706] = 'd0;
    mem[5707] = 'd0;
    mem[5708] = 'd340;
    mem[5709] = 'd0;
    mem[5710] = 'd820;
    mem[5711] = 'd0;
    mem[5712] = 'd0;
    mem[5713] = 'd0;
    mem[5714] = 'd392;
    mem[5715] = 'd0;
    mem[5716] = 'd980;
    mem[5717] = 'd0;
    mem[5718] = 'd0;
    mem[5719] = 'd0;
    mem[5720] = 'd396;
    mem[5721] = 'd0;
    mem[5722] = 'd988;
    mem[5723] = 'd0;
    mem[5724] = 'd0;
    mem[5725] = 'd0;
    mem[5726] = 'd396;
    mem[5727] = 'd0;
    mem[5728] = 'd984;
    mem[5729] = 'd0;
    mem[5730] = 'd0;
    mem[5731] = 'd0;
    mem[5732] = 'd396;
    mem[5733] = 'd0;
    mem[5734] = 'd988;
    mem[5735] = 'd0;
    mem[5736] = 'd0;
    mem[5737] = 'd0;
    mem[5738] = 'd396;
    mem[5739] = 'd0;
    mem[5740] = 'd988;
    mem[5741] = 'd0;
    mem[5742] = 'd0;
    mem[5743] = 'd0;
    mem[5744] = 'd380;
    mem[5745] = 'd0;
    mem[5746] = 'd944;
    mem[5747] = 'd0;
    mem[5748] = 'd0;
    mem[5749] = 'd0;
    mem[5750] = 'd336;
    mem[5751] = 'd0;
    mem[5752] = 'd788;
    mem[5753] = 'd0;
    mem[5754] = 'd0;
    mem[5755] = 'd0;
    mem[5756] = 'd296;
    mem[5757] = 'd0;
    mem[5758] = 'd596;
    mem[5759] = 'd0;
    mem[5760] = 'd0;
    mem[5761] = 'd0;
    mem[5762] = 'd244;
    mem[5763] = 'd0;
    mem[5764] = 'd408;
    mem[5765] = 'd0;
    mem[5766] = 'd0;
    mem[5767] = 'd0;
    mem[5768] = 'd200;
    mem[5769] = 'd0;
    mem[5770] = 'd288;
    mem[5771] = 'd0;
    mem[5772] = 'd0;
    mem[5773] = 'd0;
    mem[5774] = 'd172;
    mem[5775] = 'd0;
    mem[5776] = 'd212;
    mem[5777] = 'd0;
    mem[5778] = 'd0;
    mem[5779] = 'd0;
    mem[5780] = 'd152;
    mem[5781] = 'd0;
    mem[5782] = 'd172;
    mem[5783] = 'd0;
    mem[5784] = 'd0;
    mem[5785] = 'd0;
    mem[5786] = 'd144;
    mem[5787] = 'd0;
    mem[5788] = 'd164;
    mem[5789] = 'd0;
    mem[5790] = 'd0;
    mem[5791] = 'd0;
    mem[5792] = 'd144;
    mem[5793] = 'd0;
    mem[5794] = 'd156;
    mem[5795] = 'd0;
    mem[5796] = 'd0;
    mem[5797] = 'd0;
    mem[5798] = 'd156;
    mem[5799] = 'd0;
    mem[5800] = 'd168;
    mem[5801] = 'd0;
    mem[5802] = 'd0;
    mem[5803] = 'd0;
    mem[5804] = 'd156;
    mem[5805] = 'd0;
    mem[5806] = 'd172;
    mem[5807] = 'd0;
    mem[5808] = 'd0;
    mem[5809] = 'd0;
    mem[5810] = 'd152;
    mem[5811] = 'd0;
    mem[5812] = 'd172;
    mem[5813] = 'd0;
    mem[5814] = 'd0;
    mem[5815] = 'd0;
    mem[5816] = 'd132;
    mem[5817] = 'd0;
    mem[5818] = 'd168;
    mem[5819] = 'd0;
    mem[5820] = 'd0;
    mem[5821] = 'd0;
    mem[5822] = 'd44;
    mem[5823] = 'd0;
    mem[5824] = 'd540;
    mem[5825] = 'd0;
    mem[5826] = 'd0;
    mem[5827] = 'd0;
    mem[5828] = 'd332;
    mem[5829] = 'd0;
    mem[5830] = 'd668;
    mem[5831] = 'd0;
    mem[5832] = 'd0;
    mem[5833] = 'd0;
    mem[5834] = 'd1020;
    mem[5835] = 'd0;
    mem[5836] = 'd1020;
    mem[5837] = 'd0;
    mem[5838] = 'd0;
    mem[5839] = 'd0;
    mem[5840] = 'd1020;
    mem[5841] = 'd0;
    mem[5842] = 'd1020;
    mem[5843] = 'd0;
    mem[5844] = 'd0;
    mem[5845] = 'd0;
    mem[5846] = 'd1020;
    mem[5847] = 'd0;
    mem[5848] = 'd1020;
    mem[5849] = 'd0;
    mem[5850] = 'd0;
    mem[5851] = 'd1020;
    mem[5852] = 'd0;
    mem[5853] = 'd1020;
    mem[5854] = 'd0;
    mem[5855] = 'd0;
    mem[5856] = 'd0;
    mem[5857] = 'd1020;
    mem[5858] = 'd0;
    mem[5859] = 'd1020;
    mem[5860] = 'd0;
    mem[5861] = 'd0;
    mem[5862] = 'd0;
    mem[5863] = 'd676;
    mem[5864] = 'd0;
    mem[5865] = 'd952;
    mem[5866] = 'd0;
    mem[5867] = 'd0;
    mem[5868] = 'd0;
    mem[5869] = 'd460;
    mem[5870] = 'd0;
    mem[5871] = 'd732;
    mem[5872] = 'd0;
    mem[5873] = 'd0;
    mem[5874] = 'd0;
    mem[5875] = 'd168;
    mem[5876] = 'd0;
    mem[5877] = 'd184;
    mem[5878] = 'd0;
    mem[5879] = 'd0;
    mem[5880] = 'd0;
    mem[5881] = 'd168;
    mem[5882] = 'd0;
    mem[5883] = 'd172;
    mem[5884] = 'd0;
    mem[5885] = 'd0;
    mem[5886] = 'd0;
    mem[5887] = 'd168;
    mem[5888] = 'd0;
    mem[5889] = 'd168;
    mem[5890] = 'd0;
    mem[5891] = 'd0;
    mem[5892] = 'd0;
    mem[5893] = 'd160;
    mem[5894] = 'd0;
    mem[5895] = 'd160;
    mem[5896] = 'd0;
    mem[5897] = 'd0;
    mem[5898] = 'd0;
    mem[5899] = 'd152;
    mem[5900] = 'd0;
    mem[5901] = 'd156;
    mem[5902] = 'd0;
    mem[5903] = 'd0;
    mem[5904] = 'd0;
    mem[5905] = 'd160;
    mem[5906] = 'd0;
    mem[5907] = 'd160;
    mem[5908] = 'd0;
    mem[5909] = 'd0;
    mem[5910] = 'd0;
    mem[5911] = 'd176;
    mem[5912] = 'd0;
    mem[5913] = 'd176;
    mem[5914] = 'd0;
    mem[5915] = 'd0;
    mem[5916] = 'd0;
    mem[5917] = 'd220;
    mem[5918] = 'd0;
    mem[5919] = 'd220;
    mem[5920] = 'd0;
    mem[5921] = 'd0;
    mem[5922] = 'd0;
    mem[5923] = 'd304;
    mem[5924] = 'd0;
    mem[5925] = 'd308;
    mem[5926] = 'd0;
    mem[5927] = 'd0;
    mem[5928] = 'd0;
    mem[5929] = 'd428;
    mem[5930] = 'd0;
    mem[5931] = 'd436;
    mem[5932] = 'd0;
    mem[5933] = 'd0;
    mem[5934] = 'd0;
    mem[5935] = 'd628;
    mem[5936] = 'd0;
    mem[5937] = 'd636;
    mem[5938] = 'd0;
    mem[5939] = 'd0;
    mem[5940] = 'd0;
    mem[5941] = 'd820;
    mem[5942] = 'd0;
    mem[5943] = 'd840;
    mem[5944] = 'd0;
    mem[5945] = 'd0;
    mem[5946] = 'd0;
    mem[5947] = 'd980;
    mem[5948] = 'd0;
    mem[5949] = 'd1004;
    mem[5950] = 'd0;
    mem[5951] = 'd0;
    mem[5952] = 'd0;
    mem[5953] = 'd988;
    mem[5954] = 'd0;
    mem[5955] = 'd1020;
    mem[5956] = 'd0;
    mem[5957] = 'd0;
    mem[5958] = 'd0;
    mem[5959] = 'd984;
    mem[5960] = 'd0;
    mem[5961] = 'd1020;
    mem[5962] = 'd0;
    mem[5963] = 'd0;
    mem[5964] = 'd0;
    mem[5965] = 'd988;
    mem[5966] = 'd0;
    mem[5967] = 'd1020;
    mem[5968] = 'd0;
    mem[5969] = 'd0;
    mem[5970] = 'd0;
    mem[5971] = 'd988;
    mem[5972] = 'd0;
    mem[5973] = 'd1020;
    mem[5974] = 'd0;
    mem[5975] = 'd0;
    mem[5976] = 'd0;
    mem[5977] = 'd944;
    mem[5978] = 'd0;
    mem[5979] = 'd972;
    mem[5980] = 'd0;
    mem[5981] = 'd0;
    mem[5982] = 'd0;
    mem[5983] = 'd788;
    mem[5984] = 'd0;
    mem[5985] = 'd804;
    mem[5986] = 'd0;
    mem[5987] = 'd0;
    mem[5988] = 'd0;
    mem[5989] = 'd596;
    mem[5990] = 'd0;
    mem[5991] = 'd608;
    mem[5992] = 'd0;
    mem[5993] = 'd0;
    mem[5994] = 'd0;
    mem[5995] = 'd408;
    mem[5996] = 'd0;
    mem[5997] = 'd412;
    mem[5998] = 'd0;
    mem[5999] = 'd0;
    mem[6000] = 'd0;
    mem[6001] = 'd288;
    mem[6002] = 'd0;
    mem[6003] = 'd296;
    mem[6004] = 'd0;
    mem[6005] = 'd0;
    mem[6006] = 'd0;
    mem[6007] = 'd212;
    mem[6008] = 'd0;
    mem[6009] = 'd216;
    mem[6010] = 'd0;
    mem[6011] = 'd0;
    mem[6012] = 'd0;
    mem[6013] = 'd172;
    mem[6014] = 'd0;
    mem[6015] = 'd176;
    mem[6016] = 'd0;
    mem[6017] = 'd0;
    mem[6018] = 'd0;
    mem[6019] = 'd164;
    mem[6020] = 'd0;
    mem[6021] = 'd160;
    mem[6022] = 'd0;
    mem[6023] = 'd0;
    mem[6024] = 'd0;
    mem[6025] = 'd156;
    mem[6026] = 'd0;
    mem[6027] = 'd160;
    mem[6028] = 'd0;
    mem[6029] = 'd0;
    mem[6030] = 'd0;
    mem[6031] = 'd168;
    mem[6032] = 'd0;
    mem[6033] = 'd172;
    mem[6034] = 'd0;
    mem[6035] = 'd0;
    mem[6036] = 'd0;
    mem[6037] = 'd172;
    mem[6038] = 'd0;
    mem[6039] = 'd176;
    mem[6040] = 'd0;
    mem[6041] = 'd0;
    mem[6042] = 'd0;
    mem[6043] = 'd172;
    mem[6044] = 'd0;
    mem[6045] = 'd180;
    mem[6046] = 'd0;
    mem[6047] = 'd0;
    mem[6048] = 'd0;
    mem[6049] = 'd168;
    mem[6050] = 'd0;
    mem[6051] = 'd184;
    mem[6052] = 'd0;
    mem[6053] = 'd0;
    mem[6054] = 'd0;
    mem[6055] = 'd540;
    mem[6056] = 'd0;
    mem[6057] = 'd860;
    mem[6058] = 'd0;
    mem[6059] = 'd0;
    mem[6060] = 'd0;
    mem[6061] = 'd668;
    mem[6062] = 'd0;
    mem[6063] = 'd956;
    mem[6064] = 'd0;
    mem[6065] = 'd0;
    mem[6066] = 'd0;
    mem[6067] = 'd1020;
    mem[6068] = 'd0;
    mem[6069] = 'd1020;
    mem[6070] = 'd0;
    mem[6071] = 'd0;
    mem[6072] = 'd0;
    mem[6073] = 'd1020;
    mem[6074] = 'd0;
    mem[6075] = 'd1020;
    mem[6076] = 'd0;
    mem[6077] = 'd0;
    mem[6078] = 'd0;
    mem[6079] = 'd1020;
    mem[6080] = 'd0;
    mem[6081] = 'd1020;
    mem[6082] = 'd0;
    mem[6083] = 'd0;
    mem[6084] = 'd0;
    mem[6085] = 'd0;
    mem[6086] = 'd1020;
    mem[6087] = 'd0;
    mem[6088] = 'd1020;
    mem[6089] = 'd0;
    mem[6090] = 'd0;
    mem[6091] = 'd0;
    mem[6092] = 'd936;
    mem[6093] = 'd0;
    mem[6094] = 'd976;
    mem[6095] = 'd0;
    mem[6096] = 'd0;
    mem[6097] = 'd0;
    mem[6098] = 'd76;
    mem[6099] = 'd0;
    mem[6100] = 'd564;
    mem[6101] = 'd0;
    mem[6102] = 'd0;
    mem[6103] = 'd0;
    mem[6104] = 'd56;
    mem[6105] = 'd0;
    mem[6106] = 'd488;
    mem[6107] = 'd0;
    mem[6108] = 'd0;
    mem[6109] = 'd0;
    mem[6110] = 'd88;
    mem[6111] = 'd0;
    mem[6112] = 'd84;
    mem[6113] = 'd0;
    mem[6114] = 'd0;
    mem[6115] = 'd0;
    mem[6116] = 'd88;
    mem[6117] = 'd0;
    mem[6118] = 'd88;
    mem[6119] = 'd0;
    mem[6120] = 'd0;
    mem[6121] = 'd0;
    mem[6122] = 'd160;
    mem[6123] = 'd0;
    mem[6124] = 'd164;
    mem[6125] = 'd0;
    mem[6126] = 'd0;
    mem[6127] = 'd0;
    mem[6128] = 'd432;
    mem[6129] = 'd0;
    mem[6130] = 'd440;
    mem[6131] = 'd0;
    mem[6132] = 'd0;
    mem[6133] = 'd0;
    mem[6134] = 'd532;
    mem[6135] = 'd0;
    mem[6136] = 'd544;
    mem[6137] = 'd0;
    mem[6138] = 'd0;
    mem[6139] = 'd0;
    mem[6140] = 'd580;
    mem[6141] = 'd0;
    mem[6142] = 'd596;
    mem[6143] = 'd0;
    mem[6144] = 'd0;
    mem[6145] = 'd0;
    mem[6146] = 'd596;
    mem[6147] = 'd0;
    mem[6148] = 'd608;
    mem[6149] = 'd0;
    mem[6150] = 'd0;
    mem[6151] = 'd0;
    mem[6152] = 'd576;
    mem[6153] = 'd0;
    mem[6154] = 'd588;
    mem[6155] = 'd0;
    mem[6156] = 'd0;
    mem[6157] = 'd0;
    mem[6158] = 'd512;
    mem[6159] = 'd0;
    mem[6160] = 'd524;
    mem[6161] = 'd0;
    mem[6162] = 'd0;
    mem[6163] = 'd0;
    mem[6164] = 'd412;
    mem[6165] = 'd0;
    mem[6166] = 'd424;
    mem[6167] = 'd0;
    mem[6168] = 'd0;
    mem[6169] = 'd0;
    mem[6170] = 'd264;
    mem[6171] = 'd0;
    mem[6172] = 'd268;
    mem[6173] = 'd0;
    mem[6174] = 'd0;
    mem[6175] = 'd0;
    mem[6176] = 'd152;
    mem[6177] = 'd0;
    mem[6178] = 'd152;
    mem[6179] = 'd0;
    mem[6180] = 'd0;
    mem[6181] = 'd0;
    mem[6182] = 'd192;
    mem[6183] = 'd0;
    mem[6184] = 'd268;
    mem[6185] = 'd0;
    mem[6186] = 'd0;
    mem[6187] = 'd0;
    mem[6188] = 'd268;
    mem[6189] = 'd0;
    mem[6190] = 'd508;
    mem[6191] = 'd0;
    mem[6192] = 'd0;
    mem[6193] = 'd0;
    mem[6194] = 'd296;
    mem[6195] = 'd0;
    mem[6196] = 'd612;
    mem[6197] = 'd0;
    mem[6198] = 'd0;
    mem[6199] = 'd0;
    mem[6200] = 'd284;
    mem[6201] = 'd0;
    mem[6202] = 'd596;
    mem[6203] = 'd0;
    mem[6204] = 'd0;
    mem[6205] = 'd0;
    mem[6206] = 'd248;
    mem[6207] = 'd0;
    mem[6208] = 'd472;
    mem[6209] = 'd0;
    mem[6210] = 'd0;
    mem[6211] = 'd0;
    mem[6212] = 'd176;
    mem[6213] = 'd0;
    mem[6214] = 'd248;
    mem[6215] = 'd0;
    mem[6216] = 'd0;
    mem[6217] = 'd0;
    mem[6218] = 'd180;
    mem[6219] = 'd0;
    mem[6220] = 'd184;
    mem[6221] = 'd0;
    mem[6222] = 'd0;
    mem[6223] = 'd0;
    mem[6224] = 'd288;
    mem[6225] = 'd0;
    mem[6226] = 'd292;
    mem[6227] = 'd0;
    mem[6228] = 'd0;
    mem[6229] = 'd0;
    mem[6230] = 'd412;
    mem[6231] = 'd0;
    mem[6232] = 'd420;
    mem[6233] = 'd0;
    mem[6234] = 'd0;
    mem[6235] = 'd0;
    mem[6236] = 'd488;
    mem[6237] = 'd0;
    mem[6238] = 'd500;
    mem[6239] = 'd0;
    mem[6240] = 'd0;
    mem[6241] = 'd0;
    mem[6242] = 'd540;
    mem[6243] = 'd0;
    mem[6244] = 'd548;
    mem[6245] = 'd0;
    mem[6246] = 'd0;
    mem[6247] = 'd0;
    mem[6248] = 'd548;
    mem[6249] = 'd0;
    mem[6250] = 'd560;
    mem[6251] = 'd0;
    mem[6252] = 'd0;
    mem[6253] = 'd0;
    mem[6254] = 'd528;
    mem[6255] = 'd0;
    mem[6256] = 'd536;
    mem[6257] = 'd0;
    mem[6258] = 'd0;
    mem[6259] = 'd0;
    mem[6260] = 'd468;
    mem[6261] = 'd0;
    mem[6262] = 'd480;
    mem[6263] = 'd0;
    mem[6264] = 'd0;
    mem[6265] = 'd0;
    mem[6266] = 'd340;
    mem[6267] = 'd0;
    mem[6268] = 'd348;
    mem[6269] = 'd0;
    mem[6270] = 'd0;
    mem[6271] = 'd0;
    mem[6272] = 'd116;
    mem[6273] = 'd0;
    mem[6274] = 'd116;
    mem[6275] = 'd0;
    mem[6276] = 'd0;
    mem[6277] = 'd0;
    mem[6278] = 'd88;
    mem[6279] = 'd0;
    mem[6280] = 'd88;
    mem[6281] = 'd0;
    mem[6282] = 'd0;
    mem[6283] = 'd0;
    mem[6284] = 'd92;
    mem[6285] = 'd0;
    mem[6286] = 'd100;
    mem[6287] = 'd0;
    mem[6288] = 'd0;
    mem[6289] = 'd0;
    mem[6290] = 'd44;
    mem[6291] = 'd0;
    mem[6292] = 'd524;
    mem[6293] = 'd0;
    mem[6294] = 'd0;
    mem[6295] = 'd0;
    mem[6296] = 'd28;
    mem[6297] = 'd0;
    mem[6298] = 'd536;
    mem[6299] = 'd0;
    mem[6300] = 'd0;
    mem[6301] = 'd0;
    mem[6302] = 'd952;
    mem[6303] = 'd0;
    mem[6304] = 'd984;
    mem[6305] = 'd0;
    mem[6306] = 'd0;
    mem[6307] = 'd0;
    mem[6308] = 'd1020;
    mem[6309] = 'd0;
    mem[6310] = 'd1020;
    mem[6311] = 'd0;
    mem[6312] = 'd0;
    mem[6313] = 'd0;
    mem[6314] = 'd1020;
    mem[6315] = 'd0;
    mem[6316] = 'd1020;
    mem[6317] = 'd0;
    mem[6318] = 'd0;
    mem[6319] = 'd1020;
    mem[6320] = 'd0;
    mem[6321] = 'd1020;
    mem[6322] = 'd0;
    mem[6323] = 'd0;
    mem[6324] = 'd0;
    mem[6325] = 'd976;
    mem[6326] = 'd0;
    mem[6327] = 'd1000;
    mem[6328] = 'd0;
    mem[6329] = 'd0;
    mem[6330] = 'd0;
    mem[6331] = 'd564;
    mem[6332] = 'd0;
    mem[6333] = 'd940;
    mem[6334] = 'd0;
    mem[6335] = 'd0;
    mem[6336] = 'd0;
    mem[6337] = 'd488;
    mem[6338] = 'd0;
    mem[6339] = 'd744;
    mem[6340] = 'd0;
    mem[6341] = 'd0;
    mem[6342] = 'd0;
    mem[6343] = 'd84;
    mem[6344] = 'd0;
    mem[6345] = 'd84;
    mem[6346] = 'd0;
    mem[6347] = 'd0;
    mem[6348] = 'd0;
    mem[6349] = 'd88;
    mem[6350] = 'd0;
    mem[6351] = 'd88;
    mem[6352] = 'd0;
    mem[6353] = 'd0;
    mem[6354] = 'd0;
    mem[6355] = 'd164;
    mem[6356] = 'd0;
    mem[6357] = 'd164;
    mem[6358] = 'd0;
    mem[6359] = 'd0;
    mem[6360] = 'd0;
    mem[6361] = 'd440;
    mem[6362] = 'd0;
    mem[6363] = 'd432;
    mem[6364] = 'd0;
    mem[6365] = 'd0;
    mem[6366] = 'd0;
    mem[6367] = 'd544;
    mem[6368] = 'd0;
    mem[6369] = 'd536;
    mem[6370] = 'd0;
    mem[6371] = 'd0;
    mem[6372] = 'd0;
    mem[6373] = 'd596;
    mem[6374] = 'd0;
    mem[6375] = 'd584;
    mem[6376] = 'd0;
    mem[6377] = 'd0;
    mem[6378] = 'd0;
    mem[6379] = 'd608;
    mem[6380] = 'd0;
    mem[6381] = 'd600;
    mem[6382] = 'd0;
    mem[6383] = 'd0;
    mem[6384] = 'd0;
    mem[6385] = 'd588;
    mem[6386] = 'd0;
    mem[6387] = 'd576;
    mem[6388] = 'd0;
    mem[6389] = 'd0;
    mem[6390] = 'd0;
    mem[6391] = 'd524;
    mem[6392] = 'd0;
    mem[6393] = 'd516;
    mem[6394] = 'd0;
    mem[6395] = 'd0;
    mem[6396] = 'd0;
    mem[6397] = 'd424;
    mem[6398] = 'd0;
    mem[6399] = 'd416;
    mem[6400] = 'd0;
    mem[6401] = 'd0;
    mem[6402] = 'd0;
    mem[6403] = 'd268;
    mem[6404] = 'd0;
    mem[6405] = 'd264;
    mem[6406] = 'd0;
    mem[6407] = 'd0;
    mem[6408] = 'd0;
    mem[6409] = 'd152;
    mem[6410] = 'd0;
    mem[6411] = 'd152;
    mem[6412] = 'd0;
    mem[6413] = 'd0;
    mem[6414] = 'd0;
    mem[6415] = 'd268;
    mem[6416] = 'd0;
    mem[6417] = 'd272;
    mem[6418] = 'd0;
    mem[6419] = 'd0;
    mem[6420] = 'd0;
    mem[6421] = 'd508;
    mem[6422] = 'd0;
    mem[6423] = 'd516;
    mem[6424] = 'd0;
    mem[6425] = 'd0;
    mem[6426] = 'd0;
    mem[6427] = 'd612;
    mem[6428] = 'd0;
    mem[6429] = 'd620;
    mem[6430] = 'd0;
    mem[6431] = 'd0;
    mem[6432] = 'd0;
    mem[6433] = 'd596;
    mem[6434] = 'd0;
    mem[6435] = 'd604;
    mem[6436] = 'd0;
    mem[6437] = 'd0;
    mem[6438] = 'd0;
    mem[6439] = 'd472;
    mem[6440] = 'd0;
    mem[6441] = 'd480;
    mem[6442] = 'd0;
    mem[6443] = 'd0;
    mem[6444] = 'd0;
    mem[6445] = 'd248;
    mem[6446] = 'd0;
    mem[6447] = 'd252;
    mem[6448] = 'd0;
    mem[6449] = 'd0;
    mem[6450] = 'd0;
    mem[6451] = 'd184;
    mem[6452] = 'd0;
    mem[6453] = 'd184;
    mem[6454] = 'd0;
    mem[6455] = 'd0;
    mem[6456] = 'd0;
    mem[6457] = 'd292;
    mem[6458] = 'd0;
    mem[6459] = 'd288;
    mem[6460] = 'd0;
    mem[6461] = 'd0;
    mem[6462] = 'd0;
    mem[6463] = 'd420;
    mem[6464] = 'd0;
    mem[6465] = 'd416;
    mem[6466] = 'd0;
    mem[6467] = 'd0;
    mem[6468] = 'd0;
    mem[6469] = 'd500;
    mem[6470] = 'd0;
    mem[6471] = 'd492;
    mem[6472] = 'd0;
    mem[6473] = 'd0;
    mem[6474] = 'd0;
    mem[6475] = 'd548;
    mem[6476] = 'd0;
    mem[6477] = 'd540;
    mem[6478] = 'd0;
    mem[6479] = 'd0;
    mem[6480] = 'd0;
    mem[6481] = 'd560;
    mem[6482] = 'd0;
    mem[6483] = 'd548;
    mem[6484] = 'd0;
    mem[6485] = 'd0;
    mem[6486] = 'd0;
    mem[6487] = 'd536;
    mem[6488] = 'd0;
    mem[6489] = 'd528;
    mem[6490] = 'd0;
    mem[6491] = 'd0;
    mem[6492] = 'd0;
    mem[6493] = 'd480;
    mem[6494] = 'd0;
    mem[6495] = 'd468;
    mem[6496] = 'd0;
    mem[6497] = 'd0;
    mem[6498] = 'd0;
    mem[6499] = 'd348;
    mem[6500] = 'd0;
    mem[6501] = 'd340;
    mem[6502] = 'd0;
    mem[6503] = 'd0;
    mem[6504] = 'd0;
    mem[6505] = 'd116;
    mem[6506] = 'd0;
    mem[6507] = 'd116;
    mem[6508] = 'd0;
    mem[6509] = 'd0;
    mem[6510] = 'd0;
    mem[6511] = 'd88;
    mem[6512] = 'd0;
    mem[6513] = 'd88;
    mem[6514] = 'd0;
    mem[6515] = 'd0;
    mem[6516] = 'd0;
    mem[6517] = 'd100;
    mem[6518] = 'd0;
    mem[6519] = 'd100;
    mem[6520] = 'd0;
    mem[6521] = 'd0;
    mem[6522] = 'd0;
    mem[6523] = 'd524;
    mem[6524] = 'd0;
    mem[6525] = 'd796;
    mem[6526] = 'd0;
    mem[6527] = 'd0;
    mem[6528] = 'd0;
    mem[6529] = 'd536;
    mem[6530] = 'd0;
    mem[6531] = 'd932;
    mem[6532] = 'd0;
    mem[6533] = 'd0;
    mem[6534] = 'd0;
    mem[6535] = 'd984;
    mem[6536] = 'd0;
    mem[6537] = 'd1004;
    mem[6538] = 'd0;
    mem[6539] = 'd0;
    mem[6540] = 'd0;
    mem[6541] = 'd1020;
    mem[6542] = 'd0;
    mem[6543] = 'd1020;
    mem[6544] = 'd0;
    mem[6545] = 'd0;
    mem[6546] = 'd0;
    mem[6547] = 'd1020;
    mem[6548] = 'd0;
    mem[6549] = 'd1020;
    mem[6550] = 'd0;
    mem[6551] = 'd0;
    mem[6552] = 'd0;
    mem[6553] = 'd0;
    mem[6554] = 'd1020;
    mem[6555] = 'd0;
    mem[6556] = 'd1020;
    mem[6557] = 'd0;
    mem[6558] = 'd0;
    mem[6559] = 'd0;
    mem[6560] = 'd720;
    mem[6561] = 'd0;
    mem[6562] = 'd852;
    mem[6563] = 'd0;
    mem[6564] = 'd0;
    mem[6565] = 'd0;
    mem[6566] = 'd16;
    mem[6567] = 'd0;
    mem[6568] = 'd552;
    mem[6569] = 'd0;
    mem[6570] = 'd0;
    mem[6571] = 'd0;
    mem[6572] = 'd52;
    mem[6573] = 'd0;
    mem[6574] = 'd632;
    mem[6575] = 'd0;
    mem[6576] = 'd0;
    mem[6577] = 'd0;
    mem[6578] = 'd92;
    mem[6579] = 'd0;
    mem[6580] = 'd152;
    mem[6581] = 'd0;
    mem[6582] = 'd0;
    mem[6583] = 'd0;
    mem[6584] = 'd84;
    mem[6585] = 'd0;
    mem[6586] = 'd84;
    mem[6587] = 'd0;
    mem[6588] = 'd0;
    mem[6589] = 'd0;
    mem[6590] = 'd328;
    mem[6591] = 'd0;
    mem[6592] = 'd332;
    mem[6593] = 'd0;
    mem[6594] = 'd0;
    mem[6595] = 'd0;
    mem[6596] = 'd452;
    mem[6597] = 'd0;
    mem[6598] = 'd464;
    mem[6599] = 'd0;
    mem[6600] = 'd0;
    mem[6601] = 'd0;
    mem[6602] = 'd508;
    mem[6603] = 'd0;
    mem[6604] = 'd520;
    mem[6605] = 'd0;
    mem[6606] = 'd0;
    mem[6607] = 'd0;
    mem[6608] = 'd532;
    mem[6609] = 'd0;
    mem[6610] = 'd544;
    mem[6611] = 'd0;
    mem[6612] = 'd0;
    mem[6613] = 'd0;
    mem[6614] = 'd536;
    mem[6615] = 'd0;
    mem[6616] = 'd552;
    mem[6617] = 'd0;
    mem[6618] = 'd0;
    mem[6619] = 'd0;
    mem[6620] = 'd540;
    mem[6621] = 'd0;
    mem[6622] = 'd552;
    mem[6623] = 'd0;
    mem[6624] = 'd0;
    mem[6625] = 'd0;
    mem[6626] = 'd536;
    mem[6627] = 'd0;
    mem[6628] = 'd548;
    mem[6629] = 'd0;
    mem[6630] = 'd0;
    mem[6631] = 'd0;
    mem[6632] = 'd540;
    mem[6633] = 'd0;
    mem[6634] = 'd556;
    mem[6635] = 'd0;
    mem[6636] = 'd0;
    mem[6637] = 'd0;
    mem[6638] = 'd564;
    mem[6639] = 'd0;
    mem[6640] = 'd576;
    mem[6641] = 'd0;
    mem[6642] = 'd0;
    mem[6643] = 'd0;
    mem[6644] = 'd520;
    mem[6645] = 'd0;
    mem[6646] = 'd532;
    mem[6647] = 'd0;
    mem[6648] = 'd0;
    mem[6649] = 'd0;
    mem[6650] = 'd196;
    mem[6651] = 'd0;
    mem[6652] = 'd200;
    mem[6653] = 'd0;
    mem[6654] = 'd0;
    mem[6655] = 'd0;
    mem[6656] = 'd100;
    mem[6657] = 'd0;
    mem[6658] = 'd104;
    mem[6659] = 'd0;
    mem[6660] = 'd0;
    mem[6661] = 'd0;
    mem[6662] = 'd144;
    mem[6663] = 'd0;
    mem[6664] = 'd144;
    mem[6665] = 'd0;
    mem[6666] = 'd0;
    mem[6667] = 'd0;
    mem[6668] = 'd128;
    mem[6669] = 'd0;
    mem[6670] = 'd128;
    mem[6671] = 'd0;
    mem[6672] = 'd0;
    mem[6673] = 'd0;
    mem[6674] = 'd100;
    mem[6675] = 'd0;
    mem[6676] = 'd100;
    mem[6677] = 'd0;
    mem[6678] = 'd0;
    mem[6679] = 'd0;
    mem[6680] = 'd248;
    mem[6681] = 'd0;
    mem[6682] = 'd252;
    mem[6683] = 'd0;
    mem[6684] = 'd0;
    mem[6685] = 'd0;
    mem[6686] = 'd464;
    mem[6687] = 'd0;
    mem[6688] = 'd476;
    mem[6689] = 'd0;
    mem[6690] = 'd0;
    mem[6691] = 'd0;
    mem[6692] = 'd480;
    mem[6693] = 'd0;
    mem[6694] = 'd492;
    mem[6695] = 'd0;
    mem[6696] = 'd0;
    mem[6697] = 'd0;
    mem[6698] = 'd460;
    mem[6699] = 'd0;
    mem[6700] = 'd472;
    mem[6701] = 'd0;
    mem[6702] = 'd0;
    mem[6703] = 'd0;
    mem[6704] = 'd456;
    mem[6705] = 'd0;
    mem[6706] = 'd464;
    mem[6707] = 'd0;
    mem[6708] = 'd0;
    mem[6709] = 'd0;
    mem[6710] = 'd452;
    mem[6711] = 'd0;
    mem[6712] = 'd460;
    mem[6713] = 'd0;
    mem[6714] = 'd0;
    mem[6715] = 'd0;
    mem[6716] = 'd440;
    mem[6717] = 'd0;
    mem[6718] = 'd452;
    mem[6719] = 'd0;
    mem[6720] = 'd0;
    mem[6721] = 'd0;
    mem[6722] = 'd420;
    mem[6723] = 'd0;
    mem[6724] = 'd432;
    mem[6725] = 'd0;
    mem[6726] = 'd0;
    mem[6727] = 'd0;
    mem[6728] = 'd388;
    mem[6729] = 'd0;
    mem[6730] = 'd396;
    mem[6731] = 'd0;
    mem[6732] = 'd0;
    mem[6733] = 'd0;
    mem[6734] = 'd328;
    mem[6735] = 'd0;
    mem[6736] = 'd336;
    mem[6737] = 'd0;
    mem[6738] = 'd0;
    mem[6739] = 'd0;
    mem[6740] = 'd208;
    mem[6741] = 'd0;
    mem[6742] = 'd212;
    mem[6743] = 'd0;
    mem[6744] = 'd0;
    mem[6745] = 'd0;
    mem[6746] = 'd84;
    mem[6747] = 'd0;
    mem[6748] = 'd84;
    mem[6749] = 'd0;
    mem[6750] = 'd0;
    mem[6751] = 'd0;
    mem[6752] = 'd84;
    mem[6753] = 'd0;
    mem[6754] = 'd212;
    mem[6755] = 'd0;
    mem[6756] = 'd0;
    mem[6757] = 'd0;
    mem[6758] = 'd40;
    mem[6759] = 'd0;
    mem[6760] = 'd596;
    mem[6761] = 'd0;
    mem[6762] = 'd0;
    mem[6763] = 'd0;
    mem[6764] = 'd12;
    mem[6765] = 'd0;
    mem[6766] = 'd556;
    mem[6767] = 'd0;
    mem[6768] = 'd0;
    mem[6769] = 'd0;
    mem[6770] = 'd652;
    mem[6771] = 'd0;
    mem[6772] = 'd816;
    mem[6773] = 'd0;
    mem[6774] = 'd0;
    mem[6775] = 'd0;
    mem[6776] = 'd1020;
    mem[6777] = 'd0;
    mem[6778] = 'd1020;
    mem[6779] = 'd0;
    mem[6780] = 'd0;
    mem[6781] = 'd0;
    mem[6782] = 'd1020;
    mem[6783] = 'd0;
    mem[6784] = 'd1020;
    mem[6785] = 'd0;
    mem[6786] = 'd0;
    mem[6787] = 'd1020;
    mem[6788] = 'd0;
    mem[6789] = 'd1020;
    mem[6790] = 'd0;
    mem[6791] = 'd0;
    mem[6792] = 'd0;
    mem[6793] = 'd852;
    mem[6794] = 'd0;
    mem[6795] = 'd972;
    mem[6796] = 'd0;
    mem[6797] = 'd0;
    mem[6798] = 'd0;
    mem[6799] = 'd552;
    mem[6800] = 'd0;
    mem[6801] = 'd948;
    mem[6802] = 'd0;
    mem[6803] = 'd0;
    mem[6804] = 'd0;
    mem[6805] = 'd632;
    mem[6806] = 'd0;
    mem[6807] = 'd952;
    mem[6808] = 'd0;
    mem[6809] = 'd0;
    mem[6810] = 'd0;
    mem[6811] = 'd152;
    mem[6812] = 'd0;
    mem[6813] = 'd184;
    mem[6814] = 'd0;
    mem[6815] = 'd0;
    mem[6816] = 'd0;
    mem[6817] = 'd84;
    mem[6818] = 'd0;
    mem[6819] = 'd84;
    mem[6820] = 'd0;
    mem[6821] = 'd0;
    mem[6822] = 'd0;
    mem[6823] = 'd332;
    mem[6824] = 'd0;
    mem[6825] = 'd328;
    mem[6826] = 'd0;
    mem[6827] = 'd0;
    mem[6828] = 'd0;
    mem[6829] = 'd464;
    mem[6830] = 'd0;
    mem[6831] = 'd452;
    mem[6832] = 'd0;
    mem[6833] = 'd0;
    mem[6834] = 'd0;
    mem[6835] = 'd520;
    mem[6836] = 'd0;
    mem[6837] = 'd512;
    mem[6838] = 'd0;
    mem[6839] = 'd0;
    mem[6840] = 'd0;
    mem[6841] = 'd544;
    mem[6842] = 'd0;
    mem[6843] = 'd536;
    mem[6844] = 'd0;
    mem[6845] = 'd0;
    mem[6846] = 'd0;
    mem[6847] = 'd552;
    mem[6848] = 'd0;
    mem[6849] = 'd540;
    mem[6850] = 'd0;
    mem[6851] = 'd0;
    mem[6852] = 'd0;
    mem[6853] = 'd552;
    mem[6854] = 'd0;
    mem[6855] = 'd540;
    mem[6856] = 'd0;
    mem[6857] = 'd0;
    mem[6858] = 'd0;
    mem[6859] = 'd548;
    mem[6860] = 'd0;
    mem[6861] = 'd540;
    mem[6862] = 'd0;
    mem[6863] = 'd0;
    mem[6864] = 'd0;
    mem[6865] = 'd556;
    mem[6866] = 'd0;
    mem[6867] = 'd544;
    mem[6868] = 'd0;
    mem[6869] = 'd0;
    mem[6870] = 'd0;
    mem[6871] = 'd576;
    mem[6872] = 'd0;
    mem[6873] = 'd564;
    mem[6874] = 'd0;
    mem[6875] = 'd0;
    mem[6876] = 'd0;
    mem[6877] = 'd532;
    mem[6878] = 'd0;
    mem[6879] = 'd520;
    mem[6880] = 'd0;
    mem[6881] = 'd0;
    mem[6882] = 'd0;
    mem[6883] = 'd200;
    mem[6884] = 'd0;
    mem[6885] = 'd196;
    mem[6886] = 'd0;
    mem[6887] = 'd0;
    mem[6888] = 'd0;
    mem[6889] = 'd104;
    mem[6890] = 'd0;
    mem[6891] = 'd100;
    mem[6892] = 'd0;
    mem[6893] = 'd0;
    mem[6894] = 'd0;
    mem[6895] = 'd144;
    mem[6896] = 'd0;
    mem[6897] = 'd144;
    mem[6898] = 'd0;
    mem[6899] = 'd0;
    mem[6900] = 'd0;
    mem[6901] = 'd128;
    mem[6902] = 'd0;
    mem[6903] = 'd128;
    mem[6904] = 'd0;
    mem[6905] = 'd0;
    mem[6906] = 'd0;
    mem[6907] = 'd100;
    mem[6908] = 'd0;
    mem[6909] = 'd100;
    mem[6910] = 'd0;
    mem[6911] = 'd0;
    mem[6912] = 'd0;
    mem[6913] = 'd252;
    mem[6914] = 'd0;
    mem[6915] = 'd248;
    mem[6916] = 'd0;
    mem[6917] = 'd0;
    mem[6918] = 'd0;
    mem[6919] = 'd476;
    mem[6920] = 'd0;
    mem[6921] = 'd464;
    mem[6922] = 'd0;
    mem[6923] = 'd0;
    mem[6924] = 'd0;
    mem[6925] = 'd492;
    mem[6926] = 'd0;
    mem[6927] = 'd484;
    mem[6928] = 'd0;
    mem[6929] = 'd0;
    mem[6930] = 'd0;
    mem[6931] = 'd472;
    mem[6932] = 'd0;
    mem[6933] = 'd460;
    mem[6934] = 'd0;
    mem[6935] = 'd0;
    mem[6936] = 'd0;
    mem[6937] = 'd464;
    mem[6938] = 'd0;
    mem[6939] = 'd456;
    mem[6940] = 'd0;
    mem[6941] = 'd0;
    mem[6942] = 'd0;
    mem[6943] = 'd460;
    mem[6944] = 'd0;
    mem[6945] = 'd452;
    mem[6946] = 'd0;
    mem[6947] = 'd0;
    mem[6948] = 'd0;
    mem[6949] = 'd452;
    mem[6950] = 'd0;
    mem[6951] = 'd444;
    mem[6952] = 'd0;
    mem[6953] = 'd0;
    mem[6954] = 'd0;
    mem[6955] = 'd432;
    mem[6956] = 'd0;
    mem[6957] = 'd424;
    mem[6958] = 'd0;
    mem[6959] = 'd0;
    mem[6960] = 'd0;
    mem[6961] = 'd396;
    mem[6962] = 'd0;
    mem[6963] = 'd388;
    mem[6964] = 'd0;
    mem[6965] = 'd0;
    mem[6966] = 'd0;
    mem[6967] = 'd336;
    mem[6968] = 'd0;
    mem[6969] = 'd332;
    mem[6970] = 'd0;
    mem[6971] = 'd0;
    mem[6972] = 'd0;
    mem[6973] = 'd212;
    mem[6974] = 'd0;
    mem[6975] = 'd208;
    mem[6976] = 'd0;
    mem[6977] = 'd0;
    mem[6978] = 'd0;
    mem[6979] = 'd84;
    mem[6980] = 'd0;
    mem[6981] = 'd84;
    mem[6982] = 'd0;
    mem[6983] = 'd0;
    mem[6984] = 'd0;
    mem[6985] = 'd212;
    mem[6986] = 'd0;
    mem[6987] = 'd280;
    mem[6988] = 'd0;
    mem[6989] = 'd0;
    mem[6990] = 'd0;
    mem[6991] = 'd596;
    mem[6992] = 'd0;
    mem[6993] = 'd896;
    mem[6994] = 'd0;
    mem[6995] = 'd0;
    mem[6996] = 'd0;
    mem[6997] = 'd556;
    mem[6998] = 'd0;
    mem[6999] = 'd932;
    mem[7000] = 'd0;
    mem[7001] = 'd0;
    mem[7002] = 'd0;
    mem[7003] = 'd816;
    mem[7004] = 'd0;
    mem[7005] = 'd960;
    mem[7006] = 'd0;
    mem[7007] = 'd0;
    mem[7008] = 'd0;
    mem[7009] = 'd1020;
    mem[7010] = 'd0;
    mem[7011] = 'd1020;
    mem[7012] = 'd0;
    mem[7013] = 'd0;
    mem[7014] = 'd0;
    mem[7015] = 'd1020;
    mem[7016] = 'd0;
    mem[7017] = 'd1020;
    mem[7018] = 'd0;
    mem[7019] = 'd0;
    mem[7020] = 'd0;
    mem[7021] = 'd0;
    mem[7022] = 'd1020;
    mem[7023] = 'd0;
    mem[7024] = 'd1020;
    mem[7025] = 'd0;
    mem[7026] = 'd0;
    mem[7027] = 'd0;
    mem[7028] = 'd464;
    mem[7029] = 'd0;
    mem[7030] = 'd716;
    mem[7031] = 'd0;
    mem[7032] = 'd0;
    mem[7033] = 'd0;
    mem[7034] = 'd20;
    mem[7035] = 'd0;
    mem[7036] = 'd572;
    mem[7037] = 'd0;
    mem[7038] = 'd0;
    mem[7039] = 'd0;
    mem[7040] = 'd72;
    mem[7041] = 'd0;
    mem[7042] = 'd640;
    mem[7043] = 'd0;
    mem[7044] = 'd0;
    mem[7045] = 'd0;
    mem[7046] = 'd96;
    mem[7047] = 'd0;
    mem[7048] = 'd384;
    mem[7049] = 'd0;
    mem[7050] = 'd0;
    mem[7051] = 'd0;
    mem[7052] = 'd92;
    mem[7053] = 'd0;
    mem[7054] = 'd88;
    mem[7055] = 'd0;
    mem[7056] = 'd0;
    mem[7057] = 'd0;
    mem[7058] = 'd212;
    mem[7059] = 'd0;
    mem[7060] = 'd216;
    mem[7061] = 'd0;
    mem[7062] = 'd0;
    mem[7063] = 'd0;
    mem[7064] = 'd252;
    mem[7065] = 'd0;
    mem[7066] = 'd256;
    mem[7067] = 'd0;
    mem[7068] = 'd0;
    mem[7069] = 'd0;
    mem[7070] = 'd260;
    mem[7071] = 'd0;
    mem[7072] = 'd268;
    mem[7073] = 'd0;
    mem[7074] = 'd0;
    mem[7075] = 'd0;
    mem[7076] = 'd272;
    mem[7077] = 'd0;
    mem[7078] = 'd280;
    mem[7079] = 'd0;
    mem[7080] = 'd0;
    mem[7081] = 'd0;
    mem[7082] = 'd280;
    mem[7083] = 'd0;
    mem[7084] = 'd292;
    mem[7085] = 'd0;
    mem[7086] = 'd0;
    mem[7087] = 'd0;
    mem[7088] = 'd280;
    mem[7089] = 'd0;
    mem[7090] = 'd288;
    mem[7091] = 'd0;
    mem[7092] = 'd0;
    mem[7093] = 'd0;
    mem[7094] = 'd264;
    mem[7095] = 'd0;
    mem[7096] = 'd268;
    mem[7097] = 'd0;
    mem[7098] = 'd0;
    mem[7099] = 'd0;
    mem[7100] = 'd244;
    mem[7101] = 'd0;
    mem[7102] = 'd252;
    mem[7103] = 'd0;
    mem[7104] = 'd0;
    mem[7105] = 'd0;
    mem[7106] = 'd232;
    mem[7107] = 'd0;
    mem[7108] = 'd236;
    mem[7109] = 'd0;
    mem[7110] = 'd0;
    mem[7111] = 'd0;
    mem[7112] = 'd216;
    mem[7113] = 'd0;
    mem[7114] = 'd224;
    mem[7115] = 'd0;
    mem[7116] = 'd0;
    mem[7117] = 'd0;
    mem[7118] = 'd144;
    mem[7119] = 'd0;
    mem[7120] = 'd148;
    mem[7121] = 'd0;
    mem[7122] = 'd0;
    mem[7123] = 'd0;
    mem[7124] = 'd84;
    mem[7125] = 'd0;
    mem[7126] = 'd84;
    mem[7127] = 'd0;
    mem[7128] = 'd0;
    mem[7129] = 'd0;
    mem[7130] = 'd76;
    mem[7131] = 'd0;
    mem[7132] = 'd264;
    mem[7133] = 'd0;
    mem[7134] = 'd0;
    mem[7135] = 'd0;
    mem[7136] = 'd76;
    mem[7137] = 'd0;
    mem[7138] = 'd188;
    mem[7139] = 'd0;
    mem[7140] = 'd0;
    mem[7141] = 'd0;
    mem[7142] = 'd84;
    mem[7143] = 'd0;
    mem[7144] = 'd84;
    mem[7145] = 'd0;
    mem[7146] = 'd0;
    mem[7147] = 'd0;
    mem[7148] = 'd148;
    mem[7149] = 'd0;
    mem[7150] = 'd152;
    mem[7151] = 'd0;
    mem[7152] = 'd0;
    mem[7153] = 'd0;
    mem[7154] = 'd180;
    mem[7155] = 'd0;
    mem[7156] = 'd184;
    mem[7157] = 'd0;
    mem[7158] = 'd0;
    mem[7159] = 'd0;
    mem[7160] = 'd180;
    mem[7161] = 'd0;
    mem[7162] = 'd188;
    mem[7163] = 'd0;
    mem[7164] = 'd0;
    mem[7165] = 'd0;
    mem[7166] = 'd184;
    mem[7167] = 'd0;
    mem[7168] = 'd188;
    mem[7169] = 'd0;
    mem[7170] = 'd0;
    mem[7171] = 'd0;
    mem[7172] = 'd192;
    mem[7173] = 'd0;
    mem[7174] = 'd196;
    mem[7175] = 'd0;
    mem[7176] = 'd0;
    mem[7177] = 'd0;
    mem[7178] = 'd196;
    mem[7179] = 'd0;
    mem[7180] = 'd200;
    mem[7181] = 'd0;
    mem[7182] = 'd0;
    mem[7183] = 'd0;
    mem[7184] = 'd184;
    mem[7185] = 'd0;
    mem[7186] = 'd188;
    mem[7187] = 'd0;
    mem[7188] = 'd0;
    mem[7189] = 'd0;
    mem[7190] = 'd168;
    mem[7191] = 'd0;
    mem[7192] = 'd172;
    mem[7193] = 'd0;
    mem[7194] = 'd0;
    mem[7195] = 'd0;
    mem[7196] = 'd148;
    mem[7197] = 'd0;
    mem[7198] = 'd156;
    mem[7199] = 'd0;
    mem[7200] = 'd0;
    mem[7201] = 'd0;
    mem[7202] = 'd136;
    mem[7203] = 'd0;
    mem[7204] = 'd140;
    mem[7205] = 'd0;
    mem[7206] = 'd0;
    mem[7207] = 'd0;
    mem[7208] = 'd104;
    mem[7209] = 'd0;
    mem[7210] = 'd104;
    mem[7211] = 'd0;
    mem[7212] = 'd0;
    mem[7213] = 'd0;
    mem[7214] = 'd92;
    mem[7215] = 'd0;
    mem[7216] = 'd88;
    mem[7217] = 'd0;
    mem[7218] = 'd0;
    mem[7219] = 'd0;
    mem[7220] = 'd68;
    mem[7221] = 'd0;
    mem[7222] = 'd420;
    mem[7223] = 'd0;
    mem[7224] = 'd0;
    mem[7225] = 'd0;
    mem[7226] = 'd56;
    mem[7227] = 'd0;
    mem[7228] = 'd612;
    mem[7229] = 'd0;
    mem[7230] = 'd0;
    mem[7231] = 'd0;
    mem[7232] = 'd20;
    mem[7233] = 'd0;
    mem[7234] = 'd572;
    mem[7235] = 'd0;
    mem[7236] = 'd0;
    mem[7237] = 'd0;
    mem[7238] = 'd420;
    mem[7239] = 'd0;
    mem[7240] = 'd692;
    mem[7241] = 'd0;
    mem[7242] = 'd0;
    mem[7243] = 'd0;
    mem[7244] = 'd1020;
    mem[7245] = 'd0;
    mem[7246] = 'd1020;
    mem[7247] = 'd0;
    mem[7248] = 'd0;
    mem[7249] = 'd0;
    mem[7250] = 'd1020;
    mem[7251] = 'd0;
    mem[7252] = 'd1020;
    mem[7253] = 'd0;
    mem[7254] = 'd0;
    mem[7255] = 'd1020;
    mem[7256] = 'd0;
    mem[7257] = 'd1020;
    mem[7258] = 'd0;
    mem[7259] = 'd0;
    mem[7260] = 'd0;
    mem[7261] = 'd716;
    mem[7262] = 'd0;
    mem[7263] = 'd940;
    mem[7264] = 'd0;
    mem[7265] = 'd0;
    mem[7266] = 'd0;
    mem[7267] = 'd572;
    mem[7268] = 'd0;
    mem[7269] = 'd956;
    mem[7270] = 'd0;
    mem[7271] = 'd0;
    mem[7272] = 'd0;
    mem[7273] = 'd640;
    mem[7274] = 'd0;
    mem[7275] = 'd948;
    mem[7276] = 'd0;
    mem[7277] = 'd0;
    mem[7278] = 'd0;
    mem[7279] = 'd384;
    mem[7280] = 'd0;
    mem[7281] = 'd524;
    mem[7282] = 'd0;
    mem[7283] = 'd0;
    mem[7284] = 'd0;
    mem[7285] = 'd88;
    mem[7286] = 'd0;
    mem[7287] = 'd88;
    mem[7288] = 'd0;
    mem[7289] = 'd0;
    mem[7290] = 'd0;
    mem[7291] = 'd216;
    mem[7292] = 'd0;
    mem[7293] = 'd212;
    mem[7294] = 'd0;
    mem[7295] = 'd0;
    mem[7296] = 'd0;
    mem[7297] = 'd256;
    mem[7298] = 'd0;
    mem[7299] = 'd252;
    mem[7300] = 'd0;
    mem[7301] = 'd0;
    mem[7302] = 'd0;
    mem[7303] = 'd268;
    mem[7304] = 'd0;
    mem[7305] = 'd264;
    mem[7306] = 'd0;
    mem[7307] = 'd0;
    mem[7308] = 'd0;
    mem[7309] = 'd280;
    mem[7310] = 'd0;
    mem[7311] = 'd276;
    mem[7312] = 'd0;
    mem[7313] = 'd0;
    mem[7314] = 'd0;
    mem[7315] = 'd292;
    mem[7316] = 'd0;
    mem[7317] = 'd284;
    mem[7318] = 'd0;
    mem[7319] = 'd0;
    mem[7320] = 'd0;
    mem[7321] = 'd288;
    mem[7322] = 'd0;
    mem[7323] = 'd280;
    mem[7324] = 'd0;
    mem[7325] = 'd0;
    mem[7326] = 'd0;
    mem[7327] = 'd268;
    mem[7328] = 'd0;
    mem[7329] = 'd264;
    mem[7330] = 'd0;
    mem[7331] = 'd0;
    mem[7332] = 'd0;
    mem[7333] = 'd252;
    mem[7334] = 'd0;
    mem[7335] = 'd244;
    mem[7336] = 'd0;
    mem[7337] = 'd0;
    mem[7338] = 'd0;
    mem[7339] = 'd236;
    mem[7340] = 'd0;
    mem[7341] = 'd232;
    mem[7342] = 'd0;
    mem[7343] = 'd0;
    mem[7344] = 'd0;
    mem[7345] = 'd224;
    mem[7346] = 'd0;
    mem[7347] = 'd220;
    mem[7348] = 'd0;
    mem[7349] = 'd0;
    mem[7350] = 'd0;
    mem[7351] = 'd148;
    mem[7352] = 'd0;
    mem[7353] = 'd144;
    mem[7354] = 'd0;
    mem[7355] = 'd0;
    mem[7356] = 'd0;
    mem[7357] = 'd84;
    mem[7358] = 'd0;
    mem[7359] = 'd84;
    mem[7360] = 'd0;
    mem[7361] = 'd0;
    mem[7362] = 'd0;
    mem[7363] = 'd264;
    mem[7364] = 'd0;
    mem[7365] = 'd320;
    mem[7366] = 'd0;
    mem[7367] = 'd0;
    mem[7368] = 'd0;
    mem[7369] = 'd188;
    mem[7370] = 'd0;
    mem[7371] = 'd220;
    mem[7372] = 'd0;
    mem[7373] = 'd0;
    mem[7374] = 'd0;
    mem[7375] = 'd84;
    mem[7376] = 'd0;
    mem[7377] = 'd84;
    mem[7378] = 'd0;
    mem[7379] = 'd0;
    mem[7380] = 'd0;
    mem[7381] = 'd152;
    mem[7382] = 'd0;
    mem[7383] = 'd148;
    mem[7384] = 'd0;
    mem[7385] = 'd0;
    mem[7386] = 'd0;
    mem[7387] = 'd184;
    mem[7388] = 'd0;
    mem[7389] = 'd180;
    mem[7390] = 'd0;
    mem[7391] = 'd0;
    mem[7392] = 'd0;
    mem[7393] = 'd188;
    mem[7394] = 'd0;
    mem[7395] = 'd180;
    mem[7396] = 'd0;
    mem[7397] = 'd0;
    mem[7398] = 'd0;
    mem[7399] = 'd188;
    mem[7400] = 'd0;
    mem[7401] = 'd188;
    mem[7402] = 'd0;
    mem[7403] = 'd0;
    mem[7404] = 'd0;
    mem[7405] = 'd196;
    mem[7406] = 'd0;
    mem[7407] = 'd192;
    mem[7408] = 'd0;
    mem[7409] = 'd0;
    mem[7410] = 'd0;
    mem[7411] = 'd200;
    mem[7412] = 'd0;
    mem[7413] = 'd196;
    mem[7414] = 'd0;
    mem[7415] = 'd0;
    mem[7416] = 'd0;
    mem[7417] = 'd188;
    mem[7418] = 'd0;
    mem[7419] = 'd184;
    mem[7420] = 'd0;
    mem[7421] = 'd0;
    mem[7422] = 'd0;
    mem[7423] = 'd172;
    mem[7424] = 'd0;
    mem[7425] = 'd168;
    mem[7426] = 'd0;
    mem[7427] = 'd0;
    mem[7428] = 'd0;
    mem[7429] = 'd156;
    mem[7430] = 'd0;
    mem[7431] = 'd148;
    mem[7432] = 'd0;
    mem[7433] = 'd0;
    mem[7434] = 'd0;
    mem[7435] = 'd140;
    mem[7436] = 'd0;
    mem[7437] = 'd140;
    mem[7438] = 'd0;
    mem[7439] = 'd0;
    mem[7440] = 'd0;
    mem[7441] = 'd104;
    mem[7442] = 'd0;
    mem[7443] = 'd104;
    mem[7444] = 'd0;
    mem[7445] = 'd0;
    mem[7446] = 'd0;
    mem[7447] = 'd88;
    mem[7448] = 'd0;
    mem[7449] = 'd88;
    mem[7450] = 'd0;
    mem[7451] = 'd0;
    mem[7452] = 'd0;
    mem[7453] = 'd420;
    mem[7454] = 'd0;
    mem[7455] = 'd600;
    mem[7456] = 'd0;
    mem[7457] = 'd0;
    mem[7458] = 'd0;
    mem[7459] = 'd612;
    mem[7460] = 'd0;
    mem[7461] = 'd908;
    mem[7462] = 'd0;
    mem[7463] = 'd0;
    mem[7464] = 'd0;
    mem[7465] = 'd572;
    mem[7466] = 'd0;
    mem[7467] = 'd948;
    mem[7468] = 'd0;
    mem[7469] = 'd0;
    mem[7470] = 'd0;
    mem[7471] = 'd692;
    mem[7472] = 'd0;
    mem[7473] = 'd940;
    mem[7474] = 'd0;
    mem[7475] = 'd0;
    mem[7476] = 'd0;
    mem[7477] = 'd1020;
    mem[7478] = 'd0;
    mem[7479] = 'd1020;
    mem[7480] = 'd0;
    mem[7481] = 'd0;
    mem[7482] = 'd0;
    mem[7483] = 'd1020;
    mem[7484] = 'd0;
    mem[7485] = 'd1020;
    mem[7486] = 'd0;
    mem[7487] = 'd0;
    mem[7488] = 'd0;
    mem[7489] = 'd0;
    mem[7490] = 'd1020;
    mem[7491] = 'd0;
    mem[7492] = 'd1020;
    mem[7493] = 'd0;
    mem[7494] = 'd0;
    mem[7495] = 'd0;
    mem[7496] = 'd288;
    mem[7497] = 'd0;
    mem[7498] = 'd616;
    mem[7499] = 'd0;
    mem[7500] = 'd0;
    mem[7501] = 'd0;
    mem[7502] = 'd24;
    mem[7503] = 'd0;
    mem[7504] = 'd588;
    mem[7505] = 'd0;
    mem[7506] = 'd0;
    mem[7507] = 'd0;
    mem[7508] = 'd76;
    mem[7509] = 'd0;
    mem[7510] = 'd652;
    mem[7511] = 'd0;
    mem[7512] = 'd0;
    mem[7513] = 'd0;
    mem[7514] = 'd84;
    mem[7515] = 'd0;
    mem[7516] = 'd540;
    mem[7517] = 'd0;
    mem[7518] = 'd0;
    mem[7519] = 'd0;
    mem[7520] = 'd92;
    mem[7521] = 'd0;
    mem[7522] = 'd96;
    mem[7523] = 'd0;
    mem[7524] = 'd0;
    mem[7525] = 'd0;
    mem[7526] = 'd88;
    mem[7527] = 'd0;
    mem[7528] = 'd88;
    mem[7529] = 'd0;
    mem[7530] = 'd0;
    mem[7531] = 'd0;
    mem[7532] = 'd104;
    mem[7533] = 'd0;
    mem[7534] = 'd104;
    mem[7535] = 'd0;
    mem[7536] = 'd0;
    mem[7537] = 'd0;
    mem[7538] = 'd112;
    mem[7539] = 'd0;
    mem[7540] = 'd116;
    mem[7541] = 'd0;
    mem[7542] = 'd0;
    mem[7543] = 'd0;
    mem[7544] = 'd124;
    mem[7545] = 'd0;
    mem[7546] = 'd128;
    mem[7547] = 'd0;
    mem[7548] = 'd0;
    mem[7549] = 'd0;
    mem[7550] = 'd136;
    mem[7551] = 'd0;
    mem[7552] = 'd144;
    mem[7553] = 'd0;
    mem[7554] = 'd0;
    mem[7555] = 'd0;
    mem[7556] = 'd148;
    mem[7557] = 'd0;
    mem[7558] = 'd156;
    mem[7559] = 'd0;
    mem[7560] = 'd0;
    mem[7561] = 'd0;
    mem[7562] = 'd148;
    mem[7563] = 'd0;
    mem[7564] = 'd152;
    mem[7565] = 'd0;
    mem[7566] = 'd0;
    mem[7567] = 'd0;
    mem[7568] = 'd144;
    mem[7569] = 'd0;
    mem[7570] = 'd148;
    mem[7571] = 'd0;
    mem[7572] = 'd0;
    mem[7573] = 'd0;
    mem[7574] = 'd148;
    mem[7575] = 'd0;
    mem[7576] = 'd152;
    mem[7577] = 'd0;
    mem[7578] = 'd0;
    mem[7579] = 'd0;
    mem[7580] = 'd128;
    mem[7581] = 'd0;
    mem[7582] = 'd132;
    mem[7583] = 'd0;
    mem[7584] = 'd0;
    mem[7585] = 'd0;
    mem[7586] = 'd108;
    mem[7587] = 'd0;
    mem[7588] = 'd108;
    mem[7589] = 'd0;
    mem[7590] = 'd0;
    mem[7591] = 'd0;
    mem[7592] = 'd80;
    mem[7593] = 'd0;
    mem[7594] = 'd80;
    mem[7595] = 'd0;
    mem[7596] = 'd0;
    mem[7597] = 'd0;
    mem[7598] = 'd136;
    mem[7599] = 'd0;
    mem[7600] = 'd704;
    mem[7601] = 'd0;
    mem[7602] = 'd0;
    mem[7603] = 'd0;
    mem[7604] = 'd124;
    mem[7605] = 'd0;
    mem[7606] = 'd568;
    mem[7607] = 'd0;
    mem[7608] = 'd0;
    mem[7609] = 'd0;
    mem[7610] = 'd84;
    mem[7611] = 'd0;
    mem[7612] = 'd84;
    mem[7613] = 'd0;
    mem[7614] = 'd0;
    mem[7615] = 'd0;
    mem[7616] = 'd116;
    mem[7617] = 'd0;
    mem[7618] = 'd120;
    mem[7619] = 'd0;
    mem[7620] = 'd0;
    mem[7621] = 'd0;
    mem[7622] = 'd160;
    mem[7623] = 'd0;
    mem[7624] = 'd168;
    mem[7625] = 'd0;
    mem[7626] = 'd0;
    mem[7627] = 'd0;
    mem[7628] = 'd176;
    mem[7629] = 'd0;
    mem[7630] = 'd180;
    mem[7631] = 'd0;
    mem[7632] = 'd0;
    mem[7633] = 'd0;
    mem[7634] = 'd180;
    mem[7635] = 'd0;
    mem[7636] = 'd184;
    mem[7637] = 'd0;
    mem[7638] = 'd0;
    mem[7639] = 'd0;
    mem[7640] = 'd192;
    mem[7641] = 'd0;
    mem[7642] = 'd196;
    mem[7643] = 'd0;
    mem[7644] = 'd0;
    mem[7645] = 'd0;
    mem[7646] = 'd196;
    mem[7647] = 'd0;
    mem[7648] = 'd204;
    mem[7649] = 'd0;
    mem[7650] = 'd0;
    mem[7651] = 'd0;
    mem[7652] = 'd188;
    mem[7653] = 'd0;
    mem[7654] = 'd196;
    mem[7655] = 'd0;
    mem[7656] = 'd0;
    mem[7657] = 'd0;
    mem[7658] = 'd180;
    mem[7659] = 'd0;
    mem[7660] = 'd184;
    mem[7661] = 'd0;
    mem[7662] = 'd0;
    mem[7663] = 'd0;
    mem[7664] = 'd172;
    mem[7665] = 'd0;
    mem[7666] = 'd176;
    mem[7667] = 'd0;
    mem[7668] = 'd0;
    mem[7669] = 'd0;
    mem[7670] = 'd160;
    mem[7671] = 'd0;
    mem[7672] = 'd160;
    mem[7673] = 'd0;
    mem[7674] = 'd0;
    mem[7675] = 'd0;
    mem[7676] = 'd124;
    mem[7677] = 'd0;
    mem[7678] = 'd128;
    mem[7679] = 'd0;
    mem[7680] = 'd0;
    mem[7681] = 'd0;
    mem[7682] = 'd96;
    mem[7683] = 'd0;
    mem[7684] = 'd108;
    mem[7685] = 'd0;
    mem[7686] = 'd0;
    mem[7687] = 'd0;
    mem[7688] = 'd44;
    mem[7689] = 'd0;
    mem[7690] = 'd552;
    mem[7691] = 'd0;
    mem[7692] = 'd0;
    mem[7693] = 'd0;
    mem[7694] = 'd68;
    mem[7695] = 'd0;
    mem[7696] = 'd636;
    mem[7697] = 'd0;
    mem[7698] = 'd0;
    mem[7699] = 'd0;
    mem[7700] = 'd28;
    mem[7701] = 'd0;
    mem[7702] = 'd588;
    mem[7703] = 'd0;
    mem[7704] = 'd0;
    mem[7705] = 'd0;
    mem[7706] = 'd240;
    mem[7707] = 'd0;
    mem[7708] = 'd600;
    mem[7709] = 'd0;
    mem[7710] = 'd0;
    mem[7711] = 'd0;
    mem[7712] = 'd1020;
    mem[7713] = 'd0;
    mem[7714] = 'd1020;
    mem[7715] = 'd0;
    mem[7716] = 'd0;
    mem[7717] = 'd0;
    mem[7718] = 'd1020;
    mem[7719] = 'd0;
    mem[7720] = 'd1020;
    mem[7721] = 'd0;
    mem[7722] = 'd0;
    mem[7723] = 'd1020;
    mem[7724] = 'd0;
    mem[7725] = 'd1020;
    mem[7726] = 'd0;
    mem[7727] = 'd0;
    mem[7728] = 'd0;
    mem[7729] = 'd616;
    mem[7730] = 'd0;
    mem[7731] = 'd920;
    mem[7732] = 'd0;
    mem[7733] = 'd0;
    mem[7734] = 'd0;
    mem[7735] = 'd588;
    mem[7736] = 'd0;
    mem[7737] = 'd956;
    mem[7738] = 'd0;
    mem[7739] = 'd0;
    mem[7740] = 'd0;
    mem[7741] = 'd652;
    mem[7742] = 'd0;
    mem[7743] = 'd960;
    mem[7744] = 'd0;
    mem[7745] = 'd0;
    mem[7746] = 'd0;
    mem[7747] = 'd540;
    mem[7748] = 'd0;
    mem[7749] = 'd768;
    mem[7750] = 'd0;
    mem[7751] = 'd0;
    mem[7752] = 'd0;
    mem[7753] = 'd96;
    mem[7754] = 'd0;
    mem[7755] = 'd96;
    mem[7756] = 'd0;
    mem[7757] = 'd0;
    mem[7758] = 'd0;
    mem[7759] = 'd88;
    mem[7760] = 'd0;
    mem[7761] = 'd88;
    mem[7762] = 'd0;
    mem[7763] = 'd0;
    mem[7764] = 'd0;
    mem[7765] = 'd104;
    mem[7766] = 'd0;
    mem[7767] = 'd104;
    mem[7768] = 'd0;
    mem[7769] = 'd0;
    mem[7770] = 'd0;
    mem[7771] = 'd116;
    mem[7772] = 'd0;
    mem[7773] = 'd112;
    mem[7774] = 'd0;
    mem[7775] = 'd0;
    mem[7776] = 'd0;
    mem[7777] = 'd128;
    mem[7778] = 'd0;
    mem[7779] = 'd124;
    mem[7780] = 'd0;
    mem[7781] = 'd0;
    mem[7782] = 'd0;
    mem[7783] = 'd144;
    mem[7784] = 'd0;
    mem[7785] = 'd140;
    mem[7786] = 'd0;
    mem[7787] = 'd0;
    mem[7788] = 'd0;
    mem[7789] = 'd156;
    mem[7790] = 'd0;
    mem[7791] = 'd148;
    mem[7792] = 'd0;
    mem[7793] = 'd0;
    mem[7794] = 'd0;
    mem[7795] = 'd152;
    mem[7796] = 'd0;
    mem[7797] = 'd148;
    mem[7798] = 'd0;
    mem[7799] = 'd0;
    mem[7800] = 'd0;
    mem[7801] = 'd148;
    mem[7802] = 'd0;
    mem[7803] = 'd144;
    mem[7804] = 'd0;
    mem[7805] = 'd0;
    mem[7806] = 'd0;
    mem[7807] = 'd152;
    mem[7808] = 'd0;
    mem[7809] = 'd148;
    mem[7810] = 'd0;
    mem[7811] = 'd0;
    mem[7812] = 'd0;
    mem[7813] = 'd132;
    mem[7814] = 'd0;
    mem[7815] = 'd128;
    mem[7816] = 'd0;
    mem[7817] = 'd0;
    mem[7818] = 'd0;
    mem[7819] = 'd108;
    mem[7820] = 'd0;
    mem[7821] = 'd108;
    mem[7822] = 'd0;
    mem[7823] = 'd0;
    mem[7824] = 'd0;
    mem[7825] = 'd80;
    mem[7826] = 'd0;
    mem[7827] = 'd76;
    mem[7828] = 'd0;
    mem[7829] = 'd0;
    mem[7830] = 'd0;
    mem[7831] = 'd704;
    mem[7832] = 'd0;
    mem[7833] = 'd844;
    mem[7834] = 'd0;
    mem[7835] = 'd0;
    mem[7836] = 'd0;
    mem[7837] = 'd568;
    mem[7838] = 'd0;
    mem[7839] = 'd672;
    mem[7840] = 'd0;
    mem[7841] = 'd0;
    mem[7842] = 'd0;
    mem[7843] = 'd84;
    mem[7844] = 'd0;
    mem[7845] = 'd80;
    mem[7846] = 'd0;
    mem[7847] = 'd0;
    mem[7848] = 'd0;
    mem[7849] = 'd120;
    mem[7850] = 'd0;
    mem[7851] = 'd120;
    mem[7852] = 'd0;
    mem[7853] = 'd0;
    mem[7854] = 'd0;
    mem[7855] = 'd168;
    mem[7856] = 'd0;
    mem[7857] = 'd164;
    mem[7858] = 'd0;
    mem[7859] = 'd0;
    mem[7860] = 'd0;
    mem[7861] = 'd180;
    mem[7862] = 'd0;
    mem[7863] = 'd172;
    mem[7864] = 'd0;
    mem[7865] = 'd0;
    mem[7866] = 'd0;
    mem[7867] = 'd184;
    mem[7868] = 'd0;
    mem[7869] = 'd180;
    mem[7870] = 'd0;
    mem[7871] = 'd0;
    mem[7872] = 'd0;
    mem[7873] = 'd196;
    mem[7874] = 'd0;
    mem[7875] = 'd192;
    mem[7876] = 'd0;
    mem[7877] = 'd0;
    mem[7878] = 'd0;
    mem[7879] = 'd204;
    mem[7880] = 'd0;
    mem[7881] = 'd200;
    mem[7882] = 'd0;
    mem[7883] = 'd0;
    mem[7884] = 'd0;
    mem[7885] = 'd196;
    mem[7886] = 'd0;
    mem[7887] = 'd192;
    mem[7888] = 'd0;
    mem[7889] = 'd0;
    mem[7890] = 'd0;
    mem[7891] = 'd184;
    mem[7892] = 'd0;
    mem[7893] = 'd180;
    mem[7894] = 'd0;
    mem[7895] = 'd0;
    mem[7896] = 'd0;
    mem[7897] = 'd176;
    mem[7898] = 'd0;
    mem[7899] = 'd172;
    mem[7900] = 'd0;
    mem[7901] = 'd0;
    mem[7902] = 'd0;
    mem[7903] = 'd160;
    mem[7904] = 'd0;
    mem[7905] = 'd160;
    mem[7906] = 'd0;
    mem[7907] = 'd0;
    mem[7908] = 'd0;
    mem[7909] = 'd128;
    mem[7910] = 'd0;
    mem[7911] = 'd124;
    mem[7912] = 'd0;
    mem[7913] = 'd0;
    mem[7914] = 'd0;
    mem[7915] = 'd108;
    mem[7916] = 'd0;
    mem[7917] = 'd112;
    mem[7918] = 'd0;
    mem[7919] = 'd0;
    mem[7920] = 'd0;
    mem[7921] = 'd552;
    mem[7922] = 'd0;
    mem[7923] = 'd812;
    mem[7924] = 'd0;
    mem[7925] = 'd0;
    mem[7926] = 'd0;
    mem[7927] = 'd636;
    mem[7928] = 'd0;
    mem[7929] = 'd936;
    mem[7930] = 'd0;
    mem[7931] = 'd0;
    mem[7932] = 'd0;
    mem[7933] = 'd588;
    mem[7934] = 'd0;
    mem[7935] = 'd960;
    mem[7936] = 'd0;
    mem[7937] = 'd0;
    mem[7938] = 'd0;
    mem[7939] = 'd600;
    mem[7940] = 'd0;
    mem[7941] = 'd912;
    mem[7942] = 'd0;
    mem[7943] = 'd0;
    mem[7944] = 'd0;
    mem[7945] = 'd1020;
    mem[7946] = 'd0;
    mem[7947] = 'd1020;
    mem[7948] = 'd0;
    mem[7949] = 'd0;
    mem[7950] = 'd0;
    mem[7951] = 'd1020;
    mem[7952] = 'd0;
    mem[7953] = 'd1020;
    mem[7954] = 'd0;
    mem[7955] = 'd0;
    mem[7956] = 'd0;
    mem[7957] = 'd0;
    mem[7958] = 'd1020;
    mem[7959] = 'd0;
    mem[7960] = 'd1020;
    mem[7961] = 'd0;
    mem[7962] = 'd0;
    mem[7963] = 'd0;
    mem[7964] = 'd168;
    mem[7965] = 'd0;
    mem[7966] = 'd556;
    mem[7967] = 'd0;
    mem[7968] = 'd0;
    mem[7969] = 'd0;
    mem[7970] = 'd28;
    mem[7971] = 'd0;
    mem[7972] = 'd588;
    mem[7973] = 'd0;
    mem[7974] = 'd0;
    mem[7975] = 'd0;
    mem[7976] = 'd68;
    mem[7977] = 'd0;
    mem[7978] = 'd660;
    mem[7979] = 'd0;
    mem[7980] = 'd0;
    mem[7981] = 'd0;
    mem[7982] = 'd68;
    mem[7983] = 'd0;
    mem[7984] = 'd624;
    mem[7985] = 'd0;
    mem[7986] = 'd0;
    mem[7987] = 'd0;
    mem[7988] = 'd88;
    mem[7989] = 'd0;
    mem[7990] = 'd192;
    mem[7991] = 'd0;
    mem[7992] = 'd0;
    mem[7993] = 'd0;
    mem[7994] = 'd108;
    mem[7995] = 'd0;
    mem[7996] = 'd108;
    mem[7997] = 'd0;
    mem[7998] = 'd0;
    mem[7999] = 'd0;
    mem[8000] = 'd132;
    mem[8001] = 'd0;
    mem[8002] = 'd136;
    mem[8003] = 'd0;
    mem[8004] = 'd0;
    mem[8005] = 'd0;
    mem[8006] = 'd164;
    mem[8007] = 'd0;
    mem[8008] = 'd168;
    mem[8009] = 'd0;
    mem[8010] = 'd0;
    mem[8011] = 'd0;
    mem[8012] = 'd176;
    mem[8013] = 'd0;
    mem[8014] = 'd180;
    mem[8015] = 'd0;
    mem[8016] = 'd0;
    mem[8017] = 'd0;
    mem[8018] = 'd180;
    mem[8019] = 'd0;
    mem[8020] = 'd184;
    mem[8021] = 'd0;
    mem[8022] = 'd0;
    mem[8023] = 'd0;
    mem[8024] = 'd180;
    mem[8025] = 'd0;
    mem[8026] = 'd184;
    mem[8027] = 'd0;
    mem[8028] = 'd0;
    mem[8029] = 'd0;
    mem[8030] = 'd184;
    mem[8031] = 'd0;
    mem[8032] = 'd192;
    mem[8033] = 'd0;
    mem[8034] = 'd0;
    mem[8035] = 'd0;
    mem[8036] = 'd188;
    mem[8037] = 'd0;
    mem[8038] = 'd196;
    mem[8039] = 'd0;
    mem[8040] = 'd0;
    mem[8041] = 'd0;
    mem[8042] = 'd180;
    mem[8043] = 'd0;
    mem[8044] = 'd184;
    mem[8045] = 'd0;
    mem[8046] = 'd0;
    mem[8047] = 'd0;
    mem[8048] = 'd128;
    mem[8049] = 'd0;
    mem[8050] = 'd132;
    mem[8051] = 'd0;
    mem[8052] = 'd0;
    mem[8053] = 'd0;
    mem[8054] = 'd116;
    mem[8055] = 'd0;
    mem[8056] = 'd120;
    mem[8057] = 'd0;
    mem[8058] = 'd0;
    mem[8059] = 'd0;
    mem[8060] = 'd88;
    mem[8061] = 'd0;
    mem[8062] = 'd260;
    mem[8063] = 'd0;
    mem[8064] = 'd0;
    mem[8065] = 'd0;
    mem[8066] = 'd180;
    mem[8067] = 'd0;
    mem[8068] = 'd876;
    mem[8069] = 'd0;
    mem[8070] = 'd0;
    mem[8071] = 'd0;
    mem[8072] = 'd168;
    mem[8073] = 'd0;
    mem[8074] = 'd848;
    mem[8075] = 'd0;
    mem[8076] = 'd0;
    mem[8077] = 'd0;
    mem[8078] = 'd80;
    mem[8079] = 'd0;
    mem[8080] = 'd156;
    mem[8081] = 'd0;
    mem[8082] = 'd0;
    mem[8083] = 'd0;
    mem[8084] = 'd120;
    mem[8085] = 'd0;
    mem[8086] = 'd120;
    mem[8087] = 'd0;
    mem[8088] = 'd0;
    mem[8089] = 'd0;
    mem[8090] = 'd172;
    mem[8091] = 'd0;
    mem[8092] = 'd176;
    mem[8093] = 'd0;
    mem[8094] = 'd0;
    mem[8095] = 'd0;
    mem[8096] = 'd208;
    mem[8097] = 'd0;
    mem[8098] = 'd212;
    mem[8099] = 'd0;
    mem[8100] = 'd0;
    mem[8101] = 'd0;
    mem[8102] = 'd212;
    mem[8103] = 'd0;
    mem[8104] = 'd216;
    mem[8105] = 'd0;
    mem[8106] = 'd0;
    mem[8107] = 'd0;
    mem[8108] = 'd208;
    mem[8109] = 'd0;
    mem[8110] = 'd212;
    mem[8111] = 'd0;
    mem[8112] = 'd0;
    mem[8113] = 'd0;
    mem[8114] = 'd204;
    mem[8115] = 'd0;
    mem[8116] = 'd212;
    mem[8117] = 'd0;
    mem[8118] = 'd0;
    mem[8119] = 'd0;
    mem[8120] = 'd212;
    mem[8121] = 'd0;
    mem[8122] = 'd216;
    mem[8123] = 'd0;
    mem[8124] = 'd0;
    mem[8125] = 'd0;
    mem[8126] = 'd212;
    mem[8127] = 'd0;
    mem[8128] = 'd216;
    mem[8129] = 'd0;
    mem[8130] = 'd0;
    mem[8131] = 'd0;
    mem[8132] = 'd200;
    mem[8133] = 'd0;
    mem[8134] = 'd204;
    mem[8135] = 'd0;
    mem[8136] = 'd0;
    mem[8137] = 'd0;
    mem[8138] = 'd160;
    mem[8139] = 'd0;
    mem[8140] = 'd164;
    mem[8141] = 'd0;
    mem[8142] = 'd0;
    mem[8143] = 'd0;
    mem[8144] = 'd136;
    mem[8145] = 'd0;
    mem[8146] = 'd136;
    mem[8147] = 'd0;
    mem[8148] = 'd0;
    mem[8149] = 'd0;
    mem[8150] = 'd76;
    mem[8151] = 'd0;
    mem[8152] = 'd224;
    mem[8153] = 'd0;
    mem[8154] = 'd0;
    mem[8155] = 'd0;
    mem[8156] = 'd40;
    mem[8157] = 'd0;
    mem[8158] = 'd596;
    mem[8159] = 'd0;
    mem[8160] = 'd0;
    mem[8161] = 'd0;
    mem[8162] = 'd68;
    mem[8163] = 'd0;
    mem[8164] = 'd652;
    mem[8165] = 'd0;
    mem[8166] = 'd0;
    mem[8167] = 'd0;
    mem[8168] = 'd32;
    mem[8169] = 'd0;
    mem[8170] = 'd592;
    mem[8171] = 'd0;
    mem[8172] = 'd0;
    mem[8173] = 'd0;
    mem[8174] = 'd136;
    mem[8175] = 'd0;
    mem[8176] = 'd540;
    mem[8177] = 'd0;
    mem[8178] = 'd0;
    mem[8179] = 'd0;
    mem[8180] = 'd1020;
    mem[8181] = 'd0;
    mem[8182] = 'd1020;
    mem[8183] = 'd0;
    mem[8184] = 'd0;
    mem[8185] = 'd0;
    mem[8186] = 'd1020;
    mem[8187] = 'd0;
    mem[8188] = 'd1020;
    mem[8189] = 'd0;
    mem[8190] = 'd0;
    mem[8191] = 'd1020;
    mem[8192] = 'd0;
    mem[8193] = 'd1020;
    mem[8194] = 'd0;
    mem[8195] = 'd0;
    mem[8196] = 'd0;
    mem[8197] = 'd556;
    mem[8198] = 'd0;
    mem[8199] = 'd896;
    mem[8200] = 'd0;
    mem[8201] = 'd0;
    mem[8202] = 'd0;
    mem[8203] = 'd588;
    mem[8204] = 'd0;
    mem[8205] = 'd956;
    mem[8206] = 'd0;
    mem[8207] = 'd0;
    mem[8208] = 'd0;
    mem[8209] = 'd660;
    mem[8210] = 'd0;
    mem[8211] = 'd972;
    mem[8212] = 'd0;
    mem[8213] = 'd0;
    mem[8214] = 'd0;
    mem[8215] = 'd624;
    mem[8216] = 'd0;
    mem[8217] = 'd904;
    mem[8218] = 'd0;
    mem[8219] = 'd0;
    mem[8220] = 'd0;
    mem[8221] = 'd192;
    mem[8222] = 'd0;
    mem[8223] = 'd240;
    mem[8224] = 'd0;
    mem[8225] = 'd0;
    mem[8226] = 'd0;
    mem[8227] = 'd108;
    mem[8228] = 'd0;
    mem[8229] = 'd108;
    mem[8230] = 'd0;
    mem[8231] = 'd0;
    mem[8232] = 'd0;
    mem[8233] = 'd136;
    mem[8234] = 'd0;
    mem[8235] = 'd132;
    mem[8236] = 'd0;
    mem[8237] = 'd0;
    mem[8238] = 'd0;
    mem[8239] = 'd168;
    mem[8240] = 'd0;
    mem[8241] = 'd164;
    mem[8242] = 'd0;
    mem[8243] = 'd0;
    mem[8244] = 'd0;
    mem[8245] = 'd180;
    mem[8246] = 'd0;
    mem[8247] = 'd176;
    mem[8248] = 'd0;
    mem[8249] = 'd0;
    mem[8250] = 'd0;
    mem[8251] = 'd184;
    mem[8252] = 'd0;
    mem[8253] = 'd180;
    mem[8254] = 'd0;
    mem[8255] = 'd0;
    mem[8256] = 'd0;
    mem[8257] = 'd184;
    mem[8258] = 'd0;
    mem[8259] = 'd180;
    mem[8260] = 'd0;
    mem[8261] = 'd0;
    mem[8262] = 'd0;
    mem[8263] = 'd192;
    mem[8264] = 'd0;
    mem[8265] = 'd188;
    mem[8266] = 'd0;
    mem[8267] = 'd0;
    mem[8268] = 'd0;
    mem[8269] = 'd196;
    mem[8270] = 'd0;
    mem[8271] = 'd192;
    mem[8272] = 'd0;
    mem[8273] = 'd0;
    mem[8274] = 'd0;
    mem[8275] = 'd184;
    mem[8276] = 'd0;
    mem[8277] = 'd180;
    mem[8278] = 'd0;
    mem[8279] = 'd0;
    mem[8280] = 'd0;
    mem[8281] = 'd132;
    mem[8282] = 'd0;
    mem[8283] = 'd128;
    mem[8284] = 'd0;
    mem[8285] = 'd0;
    mem[8286] = 'd0;
    mem[8287] = 'd120;
    mem[8288] = 'd0;
    mem[8289] = 'd116;
    mem[8290] = 'd0;
    mem[8291] = 'd0;
    mem[8292] = 'd0;
    mem[8293] = 'd260;
    mem[8294] = 'd0;
    mem[8295] = 'd296;
    mem[8296] = 'd0;
    mem[8297] = 'd0;
    mem[8298] = 'd0;
    mem[8299] = 'd876;
    mem[8300] = 'd0;
    mem[8301] = 'd1004;
    mem[8302] = 'd0;
    mem[8303] = 'd0;
    mem[8304] = 'd0;
    mem[8305] = 'd848;
    mem[8306] = 'd0;
    mem[8307] = 'd980;
    mem[8308] = 'd0;
    mem[8309] = 'd0;
    mem[8310] = 'd0;
    mem[8311] = 'd156;
    mem[8312] = 'd0;
    mem[8313] = 'd176;
    mem[8314] = 'd0;
    mem[8315] = 'd0;
    mem[8316] = 'd0;
    mem[8317] = 'd120;
    mem[8318] = 'd0;
    mem[8319] = 'd120;
    mem[8320] = 'd0;
    mem[8321] = 'd0;
    mem[8322] = 'd0;
    mem[8323] = 'd176;
    mem[8324] = 'd0;
    mem[8325] = 'd172;
    mem[8326] = 'd0;
    mem[8327] = 'd0;
    mem[8328] = 'd0;
    mem[8329] = 'd212;
    mem[8330] = 'd0;
    mem[8331] = 'd208;
    mem[8332] = 'd0;
    mem[8333] = 'd0;
    mem[8334] = 'd0;
    mem[8335] = 'd216;
    mem[8336] = 'd0;
    mem[8337] = 'd212;
    mem[8338] = 'd0;
    mem[8339] = 'd0;
    mem[8340] = 'd0;
    mem[8341] = 'd212;
    mem[8342] = 'd0;
    mem[8343] = 'd208;
    mem[8344] = 'd0;
    mem[8345] = 'd0;
    mem[8346] = 'd0;
    mem[8347] = 'd212;
    mem[8348] = 'd0;
    mem[8349] = 'd204;
    mem[8350] = 'd0;
    mem[8351] = 'd0;
    mem[8352] = 'd0;
    mem[8353] = 'd216;
    mem[8354] = 'd0;
    mem[8355] = 'd212;
    mem[8356] = 'd0;
    mem[8357] = 'd0;
    mem[8358] = 'd0;
    mem[8359] = 'd216;
    mem[8360] = 'd0;
    mem[8361] = 'd216;
    mem[8362] = 'd0;
    mem[8363] = 'd0;
    mem[8364] = 'd0;
    mem[8365] = 'd204;
    mem[8366] = 'd0;
    mem[8367] = 'd200;
    mem[8368] = 'd0;
    mem[8369] = 'd0;
    mem[8370] = 'd0;
    mem[8371] = 'd164;
    mem[8372] = 'd0;
    mem[8373] = 'd160;
    mem[8374] = 'd0;
    mem[8375] = 'd0;
    mem[8376] = 'd0;
    mem[8377] = 'd136;
    mem[8378] = 'd0;
    mem[8379] = 'd136;
    mem[8380] = 'd0;
    mem[8381] = 'd0;
    mem[8382] = 'd0;
    mem[8383] = 'd224;
    mem[8384] = 'd0;
    mem[8385] = 'd304;
    mem[8386] = 'd0;
    mem[8387] = 'd0;
    mem[8388] = 'd0;
    mem[8389] = 'd596;
    mem[8390] = 'd0;
    mem[8391] = 'd880;
    mem[8392] = 'd0;
    mem[8393] = 'd0;
    mem[8394] = 'd0;
    mem[8395] = 'd652;
    mem[8396] = 'd0;
    mem[8397] = 'd960;
    mem[8398] = 'd0;
    mem[8399] = 'd0;
    mem[8400] = 'd0;
    mem[8401] = 'd592;
    mem[8402] = 'd0;
    mem[8403] = 'd956;
    mem[8404] = 'd0;
    mem[8405] = 'd0;
    mem[8406] = 'd0;
    mem[8407] = 'd540;
    mem[8408] = 'd0;
    mem[8409] = 'd892;
    mem[8410] = 'd0;
    mem[8411] = 'd0;
    mem[8412] = 'd0;
    mem[8413] = 'd1020;
    mem[8414] = 'd0;
    mem[8415] = 'd1020;
    mem[8416] = 'd0;
    mem[8417] = 'd0;
    mem[8418] = 'd0;
    mem[8419] = 'd1020;
    mem[8420] = 'd0;
    mem[8421] = 'd1020;
    mem[8422] = 'd0;
    mem[8423] = 'd0;
    mem[8424] = 'd0;
    mem[8425] = 'd0;
    mem[8426] = 'd1020;
    mem[8427] = 'd0;
    mem[8428] = 'd1020;
    mem[8429] = 'd0;
    mem[8430] = 'd0;
    mem[8431] = 'd0;
    mem[8432] = 'd124;
    mem[8433] = 'd0;
    mem[8434] = 'd528;
    mem[8435] = 'd0;
    mem[8436] = 'd0;
    mem[8437] = 'd0;
    mem[8438] = 'd28;
    mem[8439] = 'd0;
    mem[8440] = 'd584;
    mem[8441] = 'd0;
    mem[8442] = 'd0;
    mem[8443] = 'd0;
    mem[8444] = 'd60;
    mem[8445] = 'd0;
    mem[8446] = 'd664;
    mem[8447] = 'd0;
    mem[8448] = 'd0;
    mem[8449] = 'd0;
    mem[8450] = 'd72;
    mem[8451] = 'd0;
    mem[8452] = 'd648;
    mem[8453] = 'd0;
    mem[8454] = 'd0;
    mem[8455] = 'd0;
    mem[8456] = 'd76;
    mem[8457] = 'd0;
    mem[8458] = 'd408;
    mem[8459] = 'd0;
    mem[8460] = 'd0;
    mem[8461] = 'd0;
    mem[8462] = 'd120;
    mem[8463] = 'd0;
    mem[8464] = 'd120;
    mem[8465] = 'd0;
    mem[8466] = 'd0;
    mem[8467] = 'd0;
    mem[8468] = 'd120;
    mem[8469] = 'd0;
    mem[8470] = 'd124;
    mem[8471] = 'd0;
    mem[8472] = 'd0;
    mem[8473] = 'd0;
    mem[8474] = 'd168;
    mem[8475] = 'd0;
    mem[8476] = 'd168;
    mem[8477] = 'd0;
    mem[8478] = 'd0;
    mem[8479] = 'd0;
    mem[8480] = 'd188;
    mem[8481] = 'd0;
    mem[8482] = 'd188;
    mem[8483] = 'd0;
    mem[8484] = 'd0;
    mem[8485] = 'd0;
    mem[8486] = 'd192;
    mem[8487] = 'd0;
    mem[8488] = 'd192;
    mem[8489] = 'd0;
    mem[8490] = 'd0;
    mem[8491] = 'd0;
    mem[8492] = 'd192;
    mem[8493] = 'd0;
    mem[8494] = 'd196;
    mem[8495] = 'd0;
    mem[8496] = 'd0;
    mem[8497] = 'd0;
    mem[8498] = 'd192;
    mem[8499] = 'd0;
    mem[8500] = 'd200;
    mem[8501] = 'd0;
    mem[8502] = 'd0;
    mem[8503] = 'd0;
    mem[8504] = 'd188;
    mem[8505] = 'd0;
    mem[8506] = 'd188;
    mem[8507] = 'd0;
    mem[8508] = 'd0;
    mem[8509] = 'd0;
    mem[8510] = 'd140;
    mem[8511] = 'd0;
    mem[8512] = 'd144;
    mem[8513] = 'd0;
    mem[8514] = 'd0;
    mem[8515] = 'd0;
    mem[8516] = 'd124;
    mem[8517] = 'd0;
    mem[8518] = 'd124;
    mem[8519] = 'd0;
    mem[8520] = 'd0;
    mem[8521] = 'd0;
    mem[8522] = 'd88;
    mem[8523] = 'd0;
    mem[8524] = 'd84;
    mem[8525] = 'd0;
    mem[8526] = 'd0;
    mem[8527] = 'd0;
    mem[8528] = 'd136;
    mem[8529] = 'd0;
    mem[8530] = 'd644;
    mem[8531] = 'd0;
    mem[8532] = 'd0;
    mem[8533] = 'd0;
    mem[8534] = 'd192;
    mem[8535] = 'd0;
    mem[8536] = 'd888;
    mem[8537] = 'd0;
    mem[8538] = 'd0;
    mem[8539] = 'd0;
    mem[8540] = 'd188;
    mem[8541] = 'd0;
    mem[8542] = 'd880;
    mem[8543] = 'd0;
    mem[8544] = 'd0;
    mem[8545] = 'd0;
    mem[8546] = 'd120;
    mem[8547] = 'd0;
    mem[8548] = 'd540;
    mem[8549] = 'd0;
    mem[8550] = 'd0;
    mem[8551] = 'd0;
    mem[8552] = 'd100;
    mem[8553] = 'd0;
    mem[8554] = 'd96;
    mem[8555] = 'd0;
    mem[8556] = 'd0;
    mem[8557] = 'd0;
    mem[8558] = 'd128;
    mem[8559] = 'd0;
    mem[8560] = 'd132;
    mem[8561] = 'd0;
    mem[8562] = 'd0;
    mem[8563] = 'd0;
    mem[8564] = 'd176;
    mem[8565] = 'd0;
    mem[8566] = 'd180;
    mem[8567] = 'd0;
    mem[8568] = 'd0;
    mem[8569] = 'd0;
    mem[8570] = 'd204;
    mem[8571] = 'd0;
    mem[8572] = 'd208;
    mem[8573] = 'd0;
    mem[8574] = 'd0;
    mem[8575] = 'd0;
    mem[8576] = 'd204;
    mem[8577] = 'd0;
    mem[8578] = 'd208;
    mem[8579] = 'd0;
    mem[8580] = 'd0;
    mem[8581] = 'd0;
    mem[8582] = 'd200;
    mem[8583] = 'd0;
    mem[8584] = 'd208;
    mem[8585] = 'd0;
    mem[8586] = 'd0;
    mem[8587] = 'd0;
    mem[8588] = 'd204;
    mem[8589] = 'd0;
    mem[8590] = 'd208;
    mem[8591] = 'd0;
    mem[8592] = 'd0;
    mem[8593] = 'd0;
    mem[8594] = 'd204;
    mem[8595] = 'd0;
    mem[8596] = 'd208;
    mem[8597] = 'd0;
    mem[8598] = 'd0;
    mem[8599] = 'd0;
    mem[8600] = 'd176;
    mem[8601] = 'd0;
    mem[8602] = 'd180;
    mem[8603] = 'd0;
    mem[8604] = 'd0;
    mem[8605] = 'd0;
    mem[8606] = 'd116;
    mem[8607] = 'd0;
    mem[8608] = 'd120;
    mem[8609] = 'd0;
    mem[8610] = 'd0;
    mem[8611] = 'd0;
    mem[8612] = 'd120;
    mem[8613] = 'd0;
    mem[8614] = 'd116;
    mem[8615] = 'd0;
    mem[8616] = 'd0;
    mem[8617] = 'd0;
    mem[8618] = 'd48;
    mem[8619] = 'd0;
    mem[8620] = 'd444;
    mem[8621] = 'd0;
    mem[8622] = 'd0;
    mem[8623] = 'd0;
    mem[8624] = 'd56;
    mem[8625] = 'd0;
    mem[8626] = 'd620;
    mem[8627] = 'd0;
    mem[8628] = 'd0;
    mem[8629] = 'd0;
    mem[8630] = 'd64;
    mem[8631] = 'd0;
    mem[8632] = 'd664;
    mem[8633] = 'd0;
    mem[8634] = 'd0;
    mem[8635] = 'd0;
    mem[8636] = 'd28;
    mem[8637] = 'd0;
    mem[8638] = 'd588;
    mem[8639] = 'd0;
    mem[8640] = 'd0;
    mem[8641] = 'd0;
    mem[8642] = 'd88;
    mem[8643] = 'd0;
    mem[8644] = 'd512;
    mem[8645] = 'd0;
    mem[8646] = 'd0;
    mem[8647] = 'd0;
    mem[8648] = 'd1012;
    mem[8649] = 'd0;
    mem[8650] = 'd1012;
    mem[8651] = 'd0;
    mem[8652] = 'd0;
    mem[8653] = 'd0;
    mem[8654] = 'd1020;
    mem[8655] = 'd0;
    mem[8656] = 'd1020;
    mem[8657] = 'd0;
    mem[8658] = 'd0;
    mem[8659] = 'd1020;
    mem[8660] = 'd0;
    mem[8661] = 'd1020;
    mem[8662] = 'd0;
    mem[8663] = 'd0;
    mem[8664] = 'd0;
    mem[8665] = 'd528;
    mem[8666] = 'd0;
    mem[8667] = 'd880;
    mem[8668] = 'd0;
    mem[8669] = 'd0;
    mem[8670] = 'd0;
    mem[8671] = 'd584;
    mem[8672] = 'd0;
    mem[8673] = 'd948;
    mem[8674] = 'd0;
    mem[8675] = 'd0;
    mem[8676] = 'd0;
    mem[8677] = 'd664;
    mem[8678] = 'd0;
    mem[8679] = 'd980;
    mem[8680] = 'd0;
    mem[8681] = 'd0;
    mem[8682] = 'd0;
    mem[8683] = 'd648;
    mem[8684] = 'd0;
    mem[8685] = 'd940;
    mem[8686] = 'd0;
    mem[8687] = 'd0;
    mem[8688] = 'd0;
    mem[8689] = 'd408;
    mem[8690] = 'd0;
    mem[8691] = 'd572;
    mem[8692] = 'd0;
    mem[8693] = 'd0;
    mem[8694] = 'd0;
    mem[8695] = 'd120;
    mem[8696] = 'd0;
    mem[8697] = 'd120;
    mem[8698] = 'd0;
    mem[8699] = 'd0;
    mem[8700] = 'd0;
    mem[8701] = 'd124;
    mem[8702] = 'd0;
    mem[8703] = 'd120;
    mem[8704] = 'd0;
    mem[8705] = 'd0;
    mem[8706] = 'd0;
    mem[8707] = 'd168;
    mem[8708] = 'd0;
    mem[8709] = 'd168;
    mem[8710] = 'd0;
    mem[8711] = 'd0;
    mem[8712] = 'd0;
    mem[8713] = 'd188;
    mem[8714] = 'd0;
    mem[8715] = 'd188;
    mem[8716] = 'd0;
    mem[8717] = 'd0;
    mem[8718] = 'd0;
    mem[8719] = 'd192;
    mem[8720] = 'd0;
    mem[8721] = 'd192;
    mem[8722] = 'd0;
    mem[8723] = 'd0;
    mem[8724] = 'd0;
    mem[8725] = 'd196;
    mem[8726] = 'd0;
    mem[8727] = 'd192;
    mem[8728] = 'd0;
    mem[8729] = 'd0;
    mem[8730] = 'd0;
    mem[8731] = 'd200;
    mem[8732] = 'd0;
    mem[8733] = 'd196;
    mem[8734] = 'd0;
    mem[8735] = 'd0;
    mem[8736] = 'd0;
    mem[8737] = 'd188;
    mem[8738] = 'd0;
    mem[8739] = 'd188;
    mem[8740] = 'd0;
    mem[8741] = 'd0;
    mem[8742] = 'd0;
    mem[8743] = 'd144;
    mem[8744] = 'd0;
    mem[8745] = 'd140;
    mem[8746] = 'd0;
    mem[8747] = 'd0;
    mem[8748] = 'd0;
    mem[8749] = 'd124;
    mem[8750] = 'd0;
    mem[8751] = 'd124;
    mem[8752] = 'd0;
    mem[8753] = 'd0;
    mem[8754] = 'd0;
    mem[8755] = 'd84;
    mem[8756] = 'd0;
    mem[8757] = 'd84;
    mem[8758] = 'd0;
    mem[8759] = 'd0;
    mem[8760] = 'd0;
    mem[8761] = 'd644;
    mem[8762] = 'd0;
    mem[8763] = 'd752;
    mem[8764] = 'd0;
    mem[8765] = 'd0;
    mem[8766] = 'd0;
    mem[8767] = 'd888;
    mem[8768] = 'd0;
    mem[8769] = 'd1016;
    mem[8770] = 'd0;
    mem[8771] = 'd0;
    mem[8772] = 'd0;
    mem[8773] = 'd880;
    mem[8774] = 'd0;
    mem[8775] = 'd1012;
    mem[8776] = 'd0;
    mem[8777] = 'd0;
    mem[8778] = 'd0;
    mem[8779] = 'd540;
    mem[8780] = 'd0;
    mem[8781] = 'd636;
    mem[8782] = 'd0;
    mem[8783] = 'd0;
    mem[8784] = 'd0;
    mem[8785] = 'd96;
    mem[8786] = 'd0;
    mem[8787] = 'd96;
    mem[8788] = 'd0;
    mem[8789] = 'd0;
    mem[8790] = 'd0;
    mem[8791] = 'd132;
    mem[8792] = 'd0;
    mem[8793] = 'd128;
    mem[8794] = 'd0;
    mem[8795] = 'd0;
    mem[8796] = 'd0;
    mem[8797] = 'd180;
    mem[8798] = 'd0;
    mem[8799] = 'd176;
    mem[8800] = 'd0;
    mem[8801] = 'd0;
    mem[8802] = 'd0;
    mem[8803] = 'd208;
    mem[8804] = 'd0;
    mem[8805] = 'd204;
    mem[8806] = 'd0;
    mem[8807] = 'd0;
    mem[8808] = 'd0;
    mem[8809] = 'd208;
    mem[8810] = 'd0;
    mem[8811] = 'd208;
    mem[8812] = 'd0;
    mem[8813] = 'd0;
    mem[8814] = 'd0;
    mem[8815] = 'd208;
    mem[8816] = 'd0;
    mem[8817] = 'd204;
    mem[8818] = 'd0;
    mem[8819] = 'd0;
    mem[8820] = 'd0;
    mem[8821] = 'd208;
    mem[8822] = 'd0;
    mem[8823] = 'd208;
    mem[8824] = 'd0;
    mem[8825] = 'd0;
    mem[8826] = 'd0;
    mem[8827] = 'd208;
    mem[8828] = 'd0;
    mem[8829] = 'd204;
    mem[8830] = 'd0;
    mem[8831] = 'd0;
    mem[8832] = 'd0;
    mem[8833] = 'd180;
    mem[8834] = 'd0;
    mem[8835] = 'd176;
    mem[8836] = 'd0;
    mem[8837] = 'd0;
    mem[8838] = 'd0;
    mem[8839] = 'd120;
    mem[8840] = 'd0;
    mem[8841] = 'd116;
    mem[8842] = 'd0;
    mem[8843] = 'd0;
    mem[8844] = 'd0;
    mem[8845] = 'd116;
    mem[8846] = 'd0;
    mem[8847] = 'd112;
    mem[8848] = 'd0;
    mem[8849] = 'd0;
    mem[8850] = 'd0;
    mem[8851] = 'd444;
    mem[8852] = 'd0;
    mem[8853] = 'd648;
    mem[8854] = 'd0;
    mem[8855] = 'd0;
    mem[8856] = 'd0;
    mem[8857] = 'd620;
    mem[8858] = 'd0;
    mem[8859] = 'd904;
    mem[8860] = 'd0;
    mem[8861] = 'd0;
    mem[8862] = 'd0;
    mem[8863] = 'd664;
    mem[8864] = 'd0;
    mem[8865] = 'd980;
    mem[8866] = 'd0;
    mem[8867] = 'd0;
    mem[8868] = 'd0;
    mem[8869] = 'd588;
    mem[8870] = 'd0;
    mem[8871] = 'd948;
    mem[8872] = 'd0;
    mem[8873] = 'd0;
    mem[8874] = 'd0;
    mem[8875] = 'd512;
    mem[8876] = 'd0;
    mem[8877] = 'd876;
    mem[8878] = 'd0;
    mem[8879] = 'd0;
    mem[8880] = 'd0;
    mem[8881] = 'd1012;
    mem[8882] = 'd0;
    mem[8883] = 'd1016;
    mem[8884] = 'd0;
    mem[8885] = 'd0;
    mem[8886] = 'd0;
    mem[8887] = 'd1020;
    mem[8888] = 'd0;
    mem[8889] = 'd1020;
    mem[8890] = 'd0;
    mem[8891] = 'd0;
    mem[8892] = 'd0;
    mem[8893] = 'd0;
    mem[8894] = 'd1020;
    mem[8895] = 'd0;
    mem[8896] = 'd1020;
    mem[8897] = 'd0;
    mem[8898] = 'd0;
    mem[8899] = 'd0;
    mem[8900] = 'd120;
    mem[8901] = 'd0;
    mem[8902] = 'd520;
    mem[8903] = 'd0;
    mem[8904] = 'd0;
    mem[8905] = 'd0;
    mem[8906] = 'd28;
    mem[8907] = 'd0;
    mem[8908] = 'd576;
    mem[8909] = 'd0;
    mem[8910] = 'd0;
    mem[8911] = 'd0;
    mem[8912] = 'd56;
    mem[8913] = 'd0;
    mem[8914] = 'd660;
    mem[8915] = 'd0;
    mem[8916] = 'd0;
    mem[8917] = 'd0;
    mem[8918] = 'd92;
    mem[8919] = 'd0;
    mem[8920] = 'd684;
    mem[8921] = 'd0;
    mem[8922] = 'd0;
    mem[8923] = 'd0;
    mem[8924] = 'd72;
    mem[8925] = 'd0;
    mem[8926] = 'd608;
    mem[8927] = 'd0;
    mem[8928] = 'd0;
    mem[8929] = 'd0;
    mem[8930] = 'd92;
    mem[8931] = 'd0;
    mem[8932] = 'd200;
    mem[8933] = 'd0;
    mem[8934] = 'd0;
    mem[8935] = 'd0;
    mem[8936] = 'd128;
    mem[8937] = 'd0;
    mem[8938] = 'd132;
    mem[8939] = 'd0;
    mem[8940] = 'd0;
    mem[8941] = 'd0;
    mem[8942] = 'd108;
    mem[8943] = 'd0;
    mem[8944] = 'd112;
    mem[8945] = 'd0;
    mem[8946] = 'd0;
    mem[8947] = 'd0;
    mem[8948] = 'd120;
    mem[8949] = 'd0;
    mem[8950] = 'd124;
    mem[8951] = 'd0;
    mem[8952] = 'd0;
    mem[8953] = 'd0;
    mem[8954] = 'd136;
    mem[8955] = 'd0;
    mem[8956] = 'd140;
    mem[8957] = 'd0;
    mem[8958] = 'd0;
    mem[8959] = 'd0;
    mem[8960] = 'd144;
    mem[8961] = 'd0;
    mem[8962] = 'd148;
    mem[8963] = 'd0;
    mem[8964] = 'd0;
    mem[8965] = 'd0;
    mem[8966] = 'd140;
    mem[8967] = 'd0;
    mem[8968] = 'd140;
    mem[8969] = 'd0;
    mem[8970] = 'd0;
    mem[8971] = 'd0;
    mem[8972] = 'd112;
    mem[8973] = 'd0;
    mem[8974] = 'd116;
    mem[8975] = 'd0;
    mem[8976] = 'd0;
    mem[8977] = 'd0;
    mem[8978] = 'd112;
    mem[8979] = 'd0;
    mem[8980] = 'd116;
    mem[8981] = 'd0;
    mem[8982] = 'd0;
    mem[8983] = 'd0;
    mem[8984] = 'd104;
    mem[8985] = 'd0;
    mem[8986] = 'd104;
    mem[8987] = 'd0;
    mem[8988] = 'd0;
    mem[8989] = 'd0;
    mem[8990] = 'd92;
    mem[8991] = 'd0;
    mem[8992] = 'd356;
    mem[8993] = 'd0;
    mem[8994] = 'd0;
    mem[8995] = 'd0;
    mem[8996] = 'd176;
    mem[8997] = 'd0;
    mem[8998] = 'd856;
    mem[8999] = 'd0;
    mem[9000] = 'd0;
    mem[9001] = 'd0;
    mem[9002] = 'd196;
    mem[9003] = 'd0;
    mem[9004] = 'd884;
    mem[9005] = 'd0;
    mem[9006] = 'd0;
    mem[9007] = 'd0;
    mem[9008] = 'd192;
    mem[9009] = 'd0;
    mem[9010] = 'd884;
    mem[9011] = 'd0;
    mem[9012] = 'd0;
    mem[9013] = 'd0;
    mem[9014] = 'd172;
    mem[9015] = 'd0;
    mem[9016] = 'd840;
    mem[9017] = 'd0;
    mem[9018] = 'd0;
    mem[9019] = 'd0;
    mem[9020] = 'd80;
    mem[9021] = 'd0;
    mem[9022] = 'd268;
    mem[9023] = 'd0;
    mem[9024] = 'd0;
    mem[9025] = 'd0;
    mem[9026] = 'd120;
    mem[9027] = 'd0;
    mem[9028] = 'd120;
    mem[9029] = 'd0;
    mem[9030] = 'd0;
    mem[9031] = 'd0;
    mem[9032] = 'd120;
    mem[9033] = 'd0;
    mem[9034] = 'd120;
    mem[9035] = 'd0;
    mem[9036] = 'd0;
    mem[9037] = 'd0;
    mem[9038] = 'd120;
    mem[9039] = 'd0;
    mem[9040] = 'd124;
    mem[9041] = 'd0;
    mem[9042] = 'd0;
    mem[9043] = 'd0;
    mem[9044] = 'd128;
    mem[9045] = 'd0;
    mem[9046] = 'd132;
    mem[9047] = 'd0;
    mem[9048] = 'd0;
    mem[9049] = 'd0;
    mem[9050] = 'd132;
    mem[9051] = 'd0;
    mem[9052] = 'd136;
    mem[9053] = 'd0;
    mem[9054] = 'd0;
    mem[9055] = 'd0;
    mem[9056] = 'd136;
    mem[9057] = 'd0;
    mem[9058] = 'd136;
    mem[9059] = 'd0;
    mem[9060] = 'd0;
    mem[9061] = 'd0;
    mem[9062] = 'd124;
    mem[9063] = 'd0;
    mem[9064] = 'd128;
    mem[9065] = 'd0;
    mem[9066] = 'd0;
    mem[9067] = 'd0;
    mem[9068] = 'd100;
    mem[9069] = 'd0;
    mem[9070] = 'd100;
    mem[9071] = 'd0;
    mem[9072] = 'd0;
    mem[9073] = 'd0;
    mem[9074] = 'd124;
    mem[9075] = 'd0;
    mem[9076] = 'd128;
    mem[9077] = 'd0;
    mem[9078] = 'd0;
    mem[9079] = 'd0;
    mem[9080] = 'd68;
    mem[9081] = 'd0;
    mem[9082] = 'd220;
    mem[9083] = 'd0;
    mem[9084] = 'd0;
    mem[9085] = 'd0;
    mem[9086] = 'd40;
    mem[9087] = 'd0;
    mem[9088] = 'd588;
    mem[9089] = 'd0;
    mem[9090] = 'd0;
    mem[9091] = 'd0;
    mem[9092] = 'd84;
    mem[9093] = 'd0;
    mem[9094] = 'd668;
    mem[9095] = 'd0;
    mem[9096] = 'd0;
    mem[9097] = 'd0;
    mem[9098] = 'd60;
    mem[9099] = 'd0;
    mem[9100] = 'd668;
    mem[9101] = 'd0;
    mem[9102] = 'd0;
    mem[9103] = 'd0;
    mem[9104] = 'd28;
    mem[9105] = 'd0;
    mem[9106] = 'd580;
    mem[9107] = 'd0;
    mem[9108] = 'd0;
    mem[9109] = 'd0;
    mem[9110] = 'd88;
    mem[9111] = 'd0;
    mem[9112] = 'd504;
    mem[9113] = 'd0;
    mem[9114] = 'd0;
    mem[9115] = 'd0;
    mem[9116] = 'd1012;
    mem[9117] = 'd0;
    mem[9118] = 'd1012;
    mem[9119] = 'd0;
    mem[9120] = 'd0;
    mem[9121] = 'd0;
    mem[9122] = 'd1020;
    mem[9123] = 'd0;
    mem[9124] = 'd1020;
    mem[9125] = 'd0;
    mem[9126] = 'd0;
    mem[9127] = 'd1020;
    mem[9128] = 'd0;
    mem[9129] = 'd1020;
    mem[9130] = 'd0;
    mem[9131] = 'd0;
    mem[9132] = 'd0;
    mem[9133] = 'd520;
    mem[9134] = 'd0;
    mem[9135] = 'd872;
    mem[9136] = 'd0;
    mem[9137] = 'd0;
    mem[9138] = 'd0;
    mem[9139] = 'd576;
    mem[9140] = 'd0;
    mem[9141] = 'd932;
    mem[9142] = 'd0;
    mem[9143] = 'd0;
    mem[9144] = 'd0;
    mem[9145] = 'd660;
    mem[9146] = 'd0;
    mem[9147] = 'd984;
    mem[9148] = 'd0;
    mem[9149] = 'd0;
    mem[9150] = 'd0;
    mem[9151] = 'd684;
    mem[9152] = 'd0;
    mem[9153] = 'd968;
    mem[9154] = 'd0;
    mem[9155] = 'd0;
    mem[9156] = 'd0;
    mem[9157] = 'd608;
    mem[9158] = 'd0;
    mem[9159] = 'd876;
    mem[9160] = 'd0;
    mem[9161] = 'd0;
    mem[9162] = 'd0;
    mem[9163] = 'd200;
    mem[9164] = 'd0;
    mem[9165] = 'd256;
    mem[9166] = 'd0;
    mem[9167] = 'd0;
    mem[9168] = 'd0;
    mem[9169] = 'd132;
    mem[9170] = 'd0;
    mem[9171] = 'd128;
    mem[9172] = 'd0;
    mem[9173] = 'd0;
    mem[9174] = 'd0;
    mem[9175] = 'd112;
    mem[9176] = 'd0;
    mem[9177] = 'd112;
    mem[9178] = 'd0;
    mem[9179] = 'd0;
    mem[9180] = 'd0;
    mem[9181] = 'd124;
    mem[9182] = 'd0;
    mem[9183] = 'd120;
    mem[9184] = 'd0;
    mem[9185] = 'd0;
    mem[9186] = 'd0;
    mem[9187] = 'd140;
    mem[9188] = 'd0;
    mem[9189] = 'd140;
    mem[9190] = 'd0;
    mem[9191] = 'd0;
    mem[9192] = 'd0;
    mem[9193] = 'd148;
    mem[9194] = 'd0;
    mem[9195] = 'd144;
    mem[9196] = 'd0;
    mem[9197] = 'd0;
    mem[9198] = 'd0;
    mem[9199] = 'd140;
    mem[9200] = 'd0;
    mem[9201] = 'd140;
    mem[9202] = 'd0;
    mem[9203] = 'd0;
    mem[9204] = 'd0;
    mem[9205] = 'd116;
    mem[9206] = 'd0;
    mem[9207] = 'd112;
    mem[9208] = 'd0;
    mem[9209] = 'd0;
    mem[9210] = 'd0;
    mem[9211] = 'd116;
    mem[9212] = 'd0;
    mem[9213] = 'd112;
    mem[9214] = 'd0;
    mem[9215] = 'd0;
    mem[9216] = 'd0;
    mem[9217] = 'd104;
    mem[9218] = 'd0;
    mem[9219] = 'd100;
    mem[9220] = 'd0;
    mem[9221] = 'd0;
    mem[9222] = 'd0;
    mem[9223] = 'd356;
    mem[9224] = 'd0;
    mem[9225] = 'd432;
    mem[9226] = 'd0;
    mem[9227] = 'd0;
    mem[9228] = 'd0;
    mem[9229] = 'd856;
    mem[9230] = 'd0;
    mem[9231] = 'd1008;
    mem[9232] = 'd0;
    mem[9233] = 'd0;
    mem[9234] = 'd0;
    mem[9235] = 'd884;
    mem[9236] = 'd0;
    mem[9237] = 'd1020;
    mem[9238] = 'd0;
    mem[9239] = 'd0;
    mem[9240] = 'd0;
    mem[9241] = 'd884;
    mem[9242] = 'd0;
    mem[9243] = 'd1020;
    mem[9244] = 'd0;
    mem[9245] = 'd0;
    mem[9246] = 'd0;
    mem[9247] = 'd840;
    mem[9248] = 'd0;
    mem[9249] = 'd992;
    mem[9250] = 'd0;
    mem[9251] = 'd0;
    mem[9252] = 'd0;
    mem[9253] = 'd268;
    mem[9254] = 'd0;
    mem[9255] = 'd324;
    mem[9256] = 'd0;
    mem[9257] = 'd0;
    mem[9258] = 'd0;
    mem[9259] = 'd120;
    mem[9260] = 'd0;
    mem[9261] = 'd120;
    mem[9262] = 'd0;
    mem[9263] = 'd0;
    mem[9264] = 'd0;
    mem[9265] = 'd120;
    mem[9266] = 'd0;
    mem[9267] = 'd120;
    mem[9268] = 'd0;
    mem[9269] = 'd0;
    mem[9270] = 'd0;
    mem[9271] = 'd124;
    mem[9272] = 'd0;
    mem[9273] = 'd120;
    mem[9274] = 'd0;
    mem[9275] = 'd0;
    mem[9276] = 'd0;
    mem[9277] = 'd132;
    mem[9278] = 'd0;
    mem[9279] = 'd132;
    mem[9280] = 'd0;
    mem[9281] = 'd0;
    mem[9282] = 'd0;
    mem[9283] = 'd136;
    mem[9284] = 'd0;
    mem[9285] = 'd136;
    mem[9286] = 'd0;
    mem[9287] = 'd0;
    mem[9288] = 'd0;
    mem[9289] = 'd136;
    mem[9290] = 'd0;
    mem[9291] = 'd132;
    mem[9292] = 'd0;
    mem[9293] = 'd0;
    mem[9294] = 'd0;
    mem[9295] = 'd128;
    mem[9296] = 'd0;
    mem[9297] = 'd124;
    mem[9298] = 'd0;
    mem[9299] = 'd0;
    mem[9300] = 'd0;
    mem[9301] = 'd100;
    mem[9302] = 'd0;
    mem[9303] = 'd100;
    mem[9304] = 'd0;
    mem[9305] = 'd0;
    mem[9306] = 'd0;
    mem[9307] = 'd128;
    mem[9308] = 'd0;
    mem[9309] = 'd128;
    mem[9310] = 'd0;
    mem[9311] = 'd0;
    mem[9312] = 'd0;
    mem[9313] = 'd220;
    mem[9314] = 'd0;
    mem[9315] = 'd300;
    mem[9316] = 'd0;
    mem[9317] = 'd0;
    mem[9318] = 'd0;
    mem[9319] = 'd588;
    mem[9320] = 'd0;
    mem[9321] = 'd872;
    mem[9322] = 'd0;
    mem[9323] = 'd0;
    mem[9324] = 'd0;
    mem[9325] = 'd668;
    mem[9326] = 'd0;
    mem[9327] = 'd956;
    mem[9328] = 'd0;
    mem[9329] = 'd0;
    mem[9330] = 'd0;
    mem[9331] = 'd668;
    mem[9332] = 'd0;
    mem[9333] = 'd984;
    mem[9334] = 'd0;
    mem[9335] = 'd0;
    mem[9336] = 'd0;
    mem[9337] = 'd580;
    mem[9338] = 'd0;
    mem[9339] = 'd940;
    mem[9340] = 'd0;
    mem[9341] = 'd0;
    mem[9342] = 'd0;
    mem[9343] = 'd504;
    mem[9344] = 'd0;
    mem[9345] = 'd872;
    mem[9346] = 'd0;
    mem[9347] = 'd0;
    mem[9348] = 'd0;
    mem[9349] = 'd1012;
    mem[9350] = 'd0;
    mem[9351] = 'd1016;
    mem[9352] = 'd0;
    mem[9353] = 'd0;
    mem[9354] = 'd0;
    mem[9355] = 'd1020;
    mem[9356] = 'd0;
    mem[9357] = 'd1020;
    mem[9358] = 'd0;
    mem[9359] = 'd0;
    mem[9360] = 'd0;
    mem[9361] = 'd0;
    mem[9362] = 'd1020;
    mem[9363] = 'd0;
    mem[9364] = 'd1020;
    mem[9365] = 'd0;
    mem[9366] = 'd0;
    mem[9367] = 'd0;
    mem[9368] = 'd168;
    mem[9369] = 'd0;
    mem[9370] = 'd536;
    mem[9371] = 'd0;
    mem[9372] = 'd0;
    mem[9373] = 'd0;
    mem[9374] = 'd24;
    mem[9375] = 'd0;
    mem[9376] = 'd560;
    mem[9377] = 'd0;
    mem[9378] = 'd0;
    mem[9379] = 'd0;
    mem[9380] = 'd48;
    mem[9381] = 'd0;
    mem[9382] = 'd648;
    mem[9383] = 'd0;
    mem[9384] = 'd0;
    mem[9385] = 'd0;
    mem[9386] = 'd104;
    mem[9387] = 'd0;
    mem[9388] = 'd700;
    mem[9389] = 'd0;
    mem[9390] = 'd0;
    mem[9391] = 'd0;
    mem[9392] = 'd112;
    mem[9393] = 'd0;
    mem[9394] = 'd680;
    mem[9395] = 'd0;
    mem[9396] = 'd0;
    mem[9397] = 'd0;
    mem[9398] = 'd76;
    mem[9399] = 'd0;
    mem[9400] = 'd548;
    mem[9401] = 'd0;
    mem[9402] = 'd0;
    mem[9403] = 'd0;
    mem[9404] = 'd84;
    mem[9405] = 'd0;
    mem[9406] = 'd168;
    mem[9407] = 'd0;
    mem[9408] = 'd0;
    mem[9409] = 'd0;
    mem[9410] = 'd132;
    mem[9411] = 'd0;
    mem[9412] = 'd132;
    mem[9413] = 'd0;
    mem[9414] = 'd0;
    mem[9415] = 'd0;
    mem[9416] = 'd152;
    mem[9417] = 'd0;
    mem[9418] = 'd152;
    mem[9419] = 'd0;
    mem[9420] = 'd0;
    mem[9421] = 'd0;
    mem[9422] = 'd152;
    mem[9423] = 'd0;
    mem[9424] = 'd152;
    mem[9425] = 'd0;
    mem[9426] = 'd0;
    mem[9427] = 'd0;
    mem[9428] = 'd152;
    mem[9429] = 'd0;
    mem[9430] = 'd156;
    mem[9431] = 'd0;
    mem[9432] = 'd0;
    mem[9433] = 'd0;
    mem[9434] = 'd144;
    mem[9435] = 'd0;
    mem[9436] = 'd144;
    mem[9437] = 'd0;
    mem[9438] = 'd0;
    mem[9439] = 'd0;
    mem[9440] = 'd136;
    mem[9441] = 'd0;
    mem[9442] = 'd136;
    mem[9443] = 'd0;
    mem[9444] = 'd0;
    mem[9445] = 'd0;
    mem[9446] = 'd88;
    mem[9447] = 'd0;
    mem[9448] = 'd88;
    mem[9449] = 'd0;
    mem[9450] = 'd0;
    mem[9451] = 'd0;
    mem[9452] = 'd84;
    mem[9453] = 'd0;
    mem[9454] = 'd360;
    mem[9455] = 'd0;
    mem[9456] = 'd0;
    mem[9457] = 'd0;
    mem[9458] = 'd164;
    mem[9459] = 'd0;
    mem[9460] = 'd816;
    mem[9461] = 'd0;
    mem[9462] = 'd0;
    mem[9463] = 'd0;
    mem[9464] = 'd196;
    mem[9465] = 'd0;
    mem[9466] = 'd868;
    mem[9467] = 'd0;
    mem[9468] = 'd0;
    mem[9469] = 'd0;
    mem[9470] = 'd200;
    mem[9471] = 'd0;
    mem[9472] = 'd876;
    mem[9473] = 'd0;
    mem[9474] = 'd0;
    mem[9475] = 'd0;
    mem[9476] = 'd196;
    mem[9477] = 'd0;
    mem[9478] = 'd876;
    mem[9479] = 'd0;
    mem[9480] = 'd0;
    mem[9481] = 'd0;
    mem[9482] = 'd196;
    mem[9483] = 'd0;
    mem[9484] = 'd868;
    mem[9485] = 'd0;
    mem[9486] = 'd0;
    mem[9487] = 'd0;
    mem[9488] = 'd152;
    mem[9489] = 'd0;
    mem[9490] = 'd780;
    mem[9491] = 'd0;
    mem[9492] = 'd0;
    mem[9493] = 'd0;
    mem[9494] = 'd76;
    mem[9495] = 'd0;
    mem[9496] = 'd288;
    mem[9497] = 'd0;
    mem[9498] = 'd0;
    mem[9499] = 'd0;
    mem[9500] = 'd104;
    mem[9501] = 'd0;
    mem[9502] = 'd100;
    mem[9503] = 'd0;
    mem[9504] = 'd0;
    mem[9505] = 'd0;
    mem[9506] = 'd156;
    mem[9507] = 'd0;
    mem[9508] = 'd156;
    mem[9509] = 'd0;
    mem[9510] = 'd0;
    mem[9511] = 'd0;
    mem[9512] = 'd152;
    mem[9513] = 'd0;
    mem[9514] = 'd152;
    mem[9515] = 'd0;
    mem[9516] = 'd0;
    mem[9517] = 'd0;
    mem[9518] = 'd148;
    mem[9519] = 'd0;
    mem[9520] = 'd152;
    mem[9521] = 'd0;
    mem[9522] = 'd0;
    mem[9523] = 'd0;
    mem[9524] = 'd144;
    mem[9525] = 'd0;
    mem[9526] = 'd148;
    mem[9527] = 'd0;
    mem[9528] = 'd0;
    mem[9529] = 'd0;
    mem[9530] = 'd140;
    mem[9531] = 'd0;
    mem[9532] = 'd144;
    mem[9533] = 'd0;
    mem[9534] = 'd0;
    mem[9535] = 'd0;
    mem[9536] = 'd132;
    mem[9537] = 'd0;
    mem[9538] = 'd128;
    mem[9539] = 'd0;
    mem[9540] = 'd0;
    mem[9541] = 'd0;
    mem[9542] = 'd68;
    mem[9543] = 'd0;
    mem[9544] = 'd164;
    mem[9545] = 'd0;
    mem[9546] = 'd0;
    mem[9547] = 'd0;
    mem[9548] = 'd44;
    mem[9549] = 'd0;
    mem[9550] = 'd556;
    mem[9551] = 'd0;
    mem[9552] = 'd0;
    mem[9553] = 'd0;
    mem[9554] = 'd96;
    mem[9555] = 'd0;
    mem[9556] = 'd660;
    mem[9557] = 'd0;
    mem[9558] = 'd0;
    mem[9559] = 'd0;
    mem[9560] = 'd100;
    mem[9561] = 'd0;
    mem[9562] = 'd700;
    mem[9563] = 'd0;
    mem[9564] = 'd0;
    mem[9565] = 'd0;
    mem[9566] = 'd52;
    mem[9567] = 'd0;
    mem[9568] = 'd652;
    mem[9569] = 'd0;
    mem[9570] = 'd0;
    mem[9571] = 'd0;
    mem[9572] = 'd28;
    mem[9573] = 'd0;
    mem[9574] = 'd568;
    mem[9575] = 'd0;
    mem[9576] = 'd0;
    mem[9577] = 'd0;
    mem[9578] = 'd136;
    mem[9579] = 'd0;
    mem[9580] = 'd520;
    mem[9581] = 'd0;
    mem[9582] = 'd0;
    mem[9583] = 'd0;
    mem[9584] = 'd1020;
    mem[9585] = 'd0;
    mem[9586] = 'd1020;
    mem[9587] = 'd0;
    mem[9588] = 'd0;
    mem[9589] = 'd0;
    mem[9590] = 'd1020;
    mem[9591] = 'd0;
    mem[9592] = 'd1020;
    mem[9593] = 'd0;
    mem[9594] = 'd0;
    mem[9595] = 'd1020;
    mem[9596] = 'd0;
    mem[9597] = 'd1020;
    mem[9598] = 'd0;
    mem[9599] = 'd0;
    mem[9600] = 'd0;
    mem[9601] = 'd536;
    mem[9602] = 'd0;
    mem[9603] = 'd868;
    mem[9604] = 'd0;
    mem[9605] = 'd0;
    mem[9606] = 'd0;
    mem[9607] = 'd560;
    mem[9608] = 'd0;
    mem[9609] = 'd924;
    mem[9610] = 'd0;
    mem[9611] = 'd0;
    mem[9612] = 'd0;
    mem[9613] = 'd648;
    mem[9614] = 'd0;
    mem[9615] = 'd976;
    mem[9616] = 'd0;
    mem[9617] = 'd0;
    mem[9618] = 'd0;
    mem[9619] = 'd700;
    mem[9620] = 'd0;
    mem[9621] = 'd996;
    mem[9622] = 'd0;
    mem[9623] = 'd0;
    mem[9624] = 'd0;
    mem[9625] = 'd680;
    mem[9626] = 'd0;
    mem[9627] = 'd956;
    mem[9628] = 'd0;
    mem[9629] = 'd0;
    mem[9630] = 'd0;
    mem[9631] = 'd548;
    mem[9632] = 'd0;
    mem[9633] = 'd780;
    mem[9634] = 'd0;
    mem[9635] = 'd0;
    mem[9636] = 'd0;
    mem[9637] = 'd168;
    mem[9638] = 'd0;
    mem[9639] = 'd208;
    mem[9640] = 'd0;
    mem[9641] = 'd0;
    mem[9642] = 'd0;
    mem[9643] = 'd132;
    mem[9644] = 'd0;
    mem[9645] = 'd128;
    mem[9646] = 'd0;
    mem[9647] = 'd0;
    mem[9648] = 'd0;
    mem[9649] = 'd152;
    mem[9650] = 'd0;
    mem[9651] = 'd152;
    mem[9652] = 'd0;
    mem[9653] = 'd0;
    mem[9654] = 'd0;
    mem[9655] = 'd152;
    mem[9656] = 'd0;
    mem[9657] = 'd152;
    mem[9658] = 'd0;
    mem[9659] = 'd0;
    mem[9660] = 'd0;
    mem[9661] = 'd156;
    mem[9662] = 'd0;
    mem[9663] = 'd152;
    mem[9664] = 'd0;
    mem[9665] = 'd0;
    mem[9666] = 'd0;
    mem[9667] = 'd144;
    mem[9668] = 'd0;
    mem[9669] = 'd144;
    mem[9670] = 'd0;
    mem[9671] = 'd0;
    mem[9672] = 'd0;
    mem[9673] = 'd136;
    mem[9674] = 'd0;
    mem[9675] = 'd136;
    mem[9676] = 'd0;
    mem[9677] = 'd0;
    mem[9678] = 'd0;
    mem[9679] = 'd88;
    mem[9680] = 'd0;
    mem[9681] = 'd88;
    mem[9682] = 'd0;
    mem[9683] = 'd0;
    mem[9684] = 'd0;
    mem[9685] = 'd360;
    mem[9686] = 'd0;
    mem[9687] = 'd452;
    mem[9688] = 'd0;
    mem[9689] = 'd0;
    mem[9690] = 'd0;
    mem[9691] = 'd816;
    mem[9692] = 'd0;
    mem[9693] = 'd984;
    mem[9694] = 'd0;
    mem[9695] = 'd0;
    mem[9696] = 'd0;
    mem[9697] = 'd868;
    mem[9698] = 'd0;
    mem[9699] = 'd1016;
    mem[9700] = 'd0;
    mem[9701] = 'd0;
    mem[9702] = 'd0;
    mem[9703] = 'd876;
    mem[9704] = 'd0;
    mem[9705] = 'd1020;
    mem[9706] = 'd0;
    mem[9707] = 'd0;
    mem[9708] = 'd0;
    mem[9709] = 'd876;
    mem[9710] = 'd0;
    mem[9711] = 'd1020;
    mem[9712] = 'd0;
    mem[9713] = 'd0;
    mem[9714] = 'd0;
    mem[9715] = 'd868;
    mem[9716] = 'd0;
    mem[9717] = 'd1016;
    mem[9718] = 'd0;
    mem[9719] = 'd0;
    mem[9720] = 'd0;
    mem[9721] = 'd780;
    mem[9722] = 'd0;
    mem[9723] = 'd956;
    mem[9724] = 'd0;
    mem[9725] = 'd0;
    mem[9726] = 'd0;
    mem[9727] = 'd288;
    mem[9728] = 'd0;
    mem[9729] = 'd356;
    mem[9730] = 'd0;
    mem[9731] = 'd0;
    mem[9732] = 'd0;
    mem[9733] = 'd100;
    mem[9734] = 'd0;
    mem[9735] = 'd100;
    mem[9736] = 'd0;
    mem[9737] = 'd0;
    mem[9738] = 'd0;
    mem[9739] = 'd156;
    mem[9740] = 'd0;
    mem[9741] = 'd156;
    mem[9742] = 'd0;
    mem[9743] = 'd0;
    mem[9744] = 'd0;
    mem[9745] = 'd152;
    mem[9746] = 'd0;
    mem[9747] = 'd152;
    mem[9748] = 'd0;
    mem[9749] = 'd0;
    mem[9750] = 'd0;
    mem[9751] = 'd152;
    mem[9752] = 'd0;
    mem[9753] = 'd148;
    mem[9754] = 'd0;
    mem[9755] = 'd0;
    mem[9756] = 'd0;
    mem[9757] = 'd148;
    mem[9758] = 'd0;
    mem[9759] = 'd144;
    mem[9760] = 'd0;
    mem[9761] = 'd0;
    mem[9762] = 'd0;
    mem[9763] = 'd144;
    mem[9764] = 'd0;
    mem[9765] = 'd140;
    mem[9766] = 'd0;
    mem[9767] = 'd0;
    mem[9768] = 'd0;
    mem[9769] = 'd128;
    mem[9770] = 'd0;
    mem[9771] = 'd124;
    mem[9772] = 'd0;
    mem[9773] = 'd0;
    mem[9774] = 'd0;
    mem[9775] = 'd164;
    mem[9776] = 'd0;
    mem[9777] = 'd216;
    mem[9778] = 'd0;
    mem[9779] = 'd0;
    mem[9780] = 'd0;
    mem[9781] = 'd556;
    mem[9782] = 'd0;
    mem[9783] = 'd816;
    mem[9784] = 'd0;
    mem[9785] = 'd0;
    mem[9786] = 'd0;
    mem[9787] = 'd660;
    mem[9788] = 'd0;
    mem[9789] = 'd936;
    mem[9790] = 'd0;
    mem[9791] = 'd0;
    mem[9792] = 'd0;
    mem[9793] = 'd700;
    mem[9794] = 'd0;
    mem[9795] = 'd996;
    mem[9796] = 'd0;
    mem[9797] = 'd0;
    mem[9798] = 'd0;
    mem[9799] = 'd652;
    mem[9800] = 'd0;
    mem[9801] = 'd980;
    mem[9802] = 'd0;
    mem[9803] = 'd0;
    mem[9804] = 'd0;
    mem[9805] = 'd568;
    mem[9806] = 'd0;
    mem[9807] = 'd928;
    mem[9808] = 'd0;
    mem[9809] = 'd0;
    mem[9810] = 'd0;
    mem[9811] = 'd520;
    mem[9812] = 'd0;
    mem[9813] = 'd864;
    mem[9814] = 'd0;
    mem[9815] = 'd0;
    mem[9816] = 'd0;
    mem[9817] = 'd1020;
    mem[9818] = 'd0;
    mem[9819] = 'd1020;
    mem[9820] = 'd0;
    mem[9821] = 'd0;
    mem[9822] = 'd0;
    mem[9823] = 'd1020;
    mem[9824] = 'd0;
    mem[9825] = 'd1020;
    mem[9826] = 'd0;
    mem[9827] = 'd0;
    mem[9828] = 'd0;
    mem[9829] = 'd0;
    mem[9830] = 'd1020;
    mem[9831] = 'd0;
    mem[9832] = 'd1020;
    mem[9833] = 'd0;
    mem[9834] = 'd0;
    mem[9835] = 'd0;
    mem[9836] = 'd280;
    mem[9837] = 'd0;
    mem[9838] = 'd592;
    mem[9839] = 'd0;
    mem[9840] = 'd0;
    mem[9841] = 'd0;
    mem[9842] = 'd24;
    mem[9843] = 'd0;
    mem[9844] = 'd540;
    mem[9845] = 'd0;
    mem[9846] = 'd0;
    mem[9847] = 'd0;
    mem[9848] = 'd44;
    mem[9849] = 'd0;
    mem[9850] = 'd632;
    mem[9851] = 'd0;
    mem[9852] = 'd0;
    mem[9853] = 'd0;
    mem[9854] = 'd88;
    mem[9855] = 'd0;
    mem[9856] = 'd700;
    mem[9857] = 'd0;
    mem[9858] = 'd0;
    mem[9859] = 'd0;
    mem[9860] = 'd140;
    mem[9861] = 'd0;
    mem[9862] = 'd728;
    mem[9863] = 'd0;
    mem[9864] = 'd0;
    mem[9865] = 'd0;
    mem[9866] = 'd144;
    mem[9867] = 'd0;
    mem[9868] = 'd708;
    mem[9869] = 'd0;
    mem[9870] = 'd0;
    mem[9871] = 'd0;
    mem[9872] = 'd108;
    mem[9873] = 'd0;
    mem[9874] = 'd640;
    mem[9875] = 'd0;
    mem[9876] = 'd0;
    mem[9877] = 'd0;
    mem[9878] = 'd84;
    mem[9879] = 'd0;
    mem[9880] = 'd440;
    mem[9881] = 'd0;
    mem[9882] = 'd0;
    mem[9883] = 'd0;
    mem[9884] = 'd76;
    mem[9885] = 'd0;
    mem[9886] = 'd268;
    mem[9887] = 'd0;
    mem[9888] = 'd0;
    mem[9889] = 'd0;
    mem[9890] = 'd72;
    mem[9891] = 'd0;
    mem[9892] = 'd184;
    mem[9893] = 'd0;
    mem[9894] = 'd0;
    mem[9895] = 'd0;
    mem[9896] = 'd72;
    mem[9897] = 'd0;
    mem[9898] = 'd156;
    mem[9899] = 'd0;
    mem[9900] = 'd0;
    mem[9901] = 'd0;
    mem[9902] = 'd72;
    mem[9903] = 'd0;
    mem[9904] = 'd204;
    mem[9905] = 'd0;
    mem[9906] = 'd0;
    mem[9907] = 'd0;
    mem[9908] = 'd88;
    mem[9909] = 'd0;
    mem[9910] = 'd336;
    mem[9911] = 'd0;
    mem[9912] = 'd0;
    mem[9913] = 'd0;
    mem[9914] = 'd132;
    mem[9915] = 'd0;
    mem[9916] = 'd636;
    mem[9917] = 'd0;
    mem[9918] = 'd0;
    mem[9919] = 'd0;
    mem[9920] = 'd184;
    mem[9921] = 'd0;
    mem[9922] = 'd828;
    mem[9923] = 'd0;
    mem[9924] = 'd0;
    mem[9925] = 'd0;
    mem[9926] = 'd208;
    mem[9927] = 'd0;
    mem[9928] = 'd856;
    mem[9929] = 'd0;
    mem[9930] = 'd0;
    mem[9931] = 'd0;
    mem[9932] = 'd208;
    mem[9933] = 'd0;
    mem[9934] = 'd864;
    mem[9935] = 'd0;
    mem[9936] = 'd0;
    mem[9937] = 'd0;
    mem[9938] = 'd204;
    mem[9939] = 'd0;
    mem[9940] = 'd864;
    mem[9941] = 'd0;
    mem[9942] = 'd0;
    mem[9943] = 'd0;
    mem[9944] = 'd208;
    mem[9945] = 'd0;
    mem[9946] = 'd864;
    mem[9947] = 'd0;
    mem[9948] = 'd0;
    mem[9949] = 'd0;
    mem[9950] = 'd208;
    mem[9951] = 'd0;
    mem[9952] = 'd864;
    mem[9953] = 'd0;
    mem[9954] = 'd0;
    mem[9955] = 'd0;
    mem[9956] = 'd204;
    mem[9957] = 'd0;
    mem[9958] = 'd856;
    mem[9959] = 'd0;
    mem[9960] = 'd0;
    mem[9961] = 'd0;
    mem[9962] = 'd176;
    mem[9963] = 'd0;
    mem[9964] = 'd812;
    mem[9965] = 'd0;
    mem[9966] = 'd0;
    mem[9967] = 'd0;
    mem[9968] = 'd108;
    mem[9969] = 'd0;
    mem[9970] = 'd572;
    mem[9971] = 'd0;
    mem[9972] = 'd0;
    mem[9973] = 'd0;
    mem[9974] = 'd72;
    mem[9975] = 'd0;
    mem[9976] = 'd292;
    mem[9977] = 'd0;
    mem[9978] = 'd0;
    mem[9979] = 'd0;
    mem[9980] = 'd64;
    mem[9981] = 'd0;
    mem[9982] = 'd188;
    mem[9983] = 'd0;
    mem[9984] = 'd0;
    mem[9985] = 'd0;
    mem[9986] = 'd64;
    mem[9987] = 'd0;
    mem[9988] = 'd148;
    mem[9989] = 'd0;
    mem[9990] = 'd0;
    mem[9991] = 'd0;
    mem[9992] = 'd64;
    mem[9993] = 'd0;
    mem[9994] = 'd176;
    mem[9995] = 'd0;
    mem[9996] = 'd0;
    mem[9997] = 'd0;
    mem[9998] = 'd60;
    mem[9999] = 'd0;
    mem[10000] = 'd276;
    mem[10001] = 'd0;
    mem[10002] = 'd0;
    mem[10003] = 'd0;
    mem[10004] = 'd60;
    mem[10005] = 'd0;
    mem[10006] = 'd428;
    mem[10007] = 'd0;
    mem[10008] = 'd0;
    mem[10009] = 'd0;
    mem[10010] = 'd76;
    mem[10011] = 'd0;
    mem[10012] = 'd632;
    mem[10013] = 'd0;
    mem[10014] = 'd0;
    mem[10015] = 'd0;
    mem[10016] = 'd132;
    mem[10017] = 'd0;
    mem[10018] = 'd692;
    mem[10019] = 'd0;
    mem[10020] = 'd0;
    mem[10021] = 'd0;
    mem[10022] = 'd140;
    mem[10023] = 'd0;
    mem[10024] = 'd724;
    mem[10025] = 'd0;
    mem[10026] = 'd0;
    mem[10027] = 'd0;
    mem[10028] = 'd84;
    mem[10029] = 'd0;
    mem[10030] = 'd700;
    mem[10031] = 'd0;
    mem[10032] = 'd0;
    mem[10033] = 'd0;
    mem[10034] = 'd48;
    mem[10035] = 'd0;
    mem[10036] = 'd636;
    mem[10037] = 'd0;
    mem[10038] = 'd0;
    mem[10039] = 'd0;
    mem[10040] = 'd28;
    mem[10041] = 'd0;
    mem[10042] = 'd548;
    mem[10043] = 'd0;
    mem[10044] = 'd0;
    mem[10045] = 'd0;
    mem[10046] = 'd236;
    mem[10047] = 'd0;
    mem[10048] = 'd568;
    mem[10049] = 'd0;
    mem[10050] = 'd0;
    mem[10051] = 'd0;
    mem[10052] = 'd1020;
    mem[10053] = 'd0;
    mem[10054] = 'd1020;
    mem[10055] = 'd0;
    mem[10056] = 'd0;
    mem[10057] = 'd0;
    mem[10058] = 'd1020;
    mem[10059] = 'd0;
    mem[10060] = 'd1020;
    mem[10061] = 'd0;
    mem[10062] = 'd0;
    mem[10063] = 'd1020;
    mem[10064] = 'd0;
    mem[10065] = 'd1020;
    mem[10066] = 'd0;
    mem[10067] = 'd0;
    mem[10068] = 'd0;
    mem[10069] = 'd592;
    mem[10070] = 'd0;
    mem[10071] = 'd876;
    mem[10072] = 'd0;
    mem[10073] = 'd0;
    mem[10074] = 'd0;
    mem[10075] = 'd540;
    mem[10076] = 'd0;
    mem[10077] = 'd908;
    mem[10078] = 'd0;
    mem[10079] = 'd0;
    mem[10080] = 'd0;
    mem[10081] = 'd632;
    mem[10082] = 'd0;
    mem[10083] = 'd960;
    mem[10084] = 'd0;
    mem[10085] = 'd0;
    mem[10086] = 'd0;
    mem[10087] = 'd700;
    mem[10088] = 'd0;
    mem[10089] = 'd1000;
    mem[10090] = 'd0;
    mem[10091] = 'd0;
    mem[10092] = 'd0;
    mem[10093] = 'd728;
    mem[10094] = 'd0;
    mem[10095] = 'd1004;
    mem[10096] = 'd0;
    mem[10097] = 'd0;
    mem[10098] = 'd0;
    mem[10099] = 'd708;
    mem[10100] = 'd0;
    mem[10101] = 'd976;
    mem[10102] = 'd0;
    mem[10103] = 'd0;
    mem[10104] = 'd0;
    mem[10105] = 'd640;
    mem[10106] = 'd0;
    mem[10107] = 'd888;
    mem[10108] = 'd0;
    mem[10109] = 'd0;
    mem[10110] = 'd0;
    mem[10111] = 'd440;
    mem[10112] = 'd0;
    mem[10113] = 'd604;
    mem[10114] = 'd0;
    mem[10115] = 'd0;
    mem[10116] = 'd0;
    mem[10117] = 'd268;
    mem[10118] = 'd0;
    mem[10119] = 'd360;
    mem[10120] = 'd0;
    mem[10121] = 'd0;
    mem[10122] = 'd0;
    mem[10123] = 'd184;
    mem[10124] = 'd0;
    mem[10125] = 'd228;
    mem[10126] = 'd0;
    mem[10127] = 'd0;
    mem[10128] = 'd0;
    mem[10129] = 'd156;
    mem[10130] = 'd0;
    mem[10131] = 'd192;
    mem[10132] = 'd0;
    mem[10133] = 'd0;
    mem[10134] = 'd0;
    mem[10135] = 'd204;
    mem[10136] = 'd0;
    mem[10137] = 'd260;
    mem[10138] = 'd0;
    mem[10139] = 'd0;
    mem[10140] = 'd0;
    mem[10141] = 'd336;
    mem[10142] = 'd0;
    mem[10143] = 'd432;
    mem[10144] = 'd0;
    mem[10145] = 'd0;
    mem[10146] = 'd0;
    mem[10147] = 'd636;
    mem[10148] = 'd0;
    mem[10149] = 'd804;
    mem[10150] = 'd0;
    mem[10151] = 'd0;
    mem[10152] = 'd0;
    mem[10153] = 'd828;
    mem[10154] = 'd0;
    mem[10155] = 'd1004;
    mem[10156] = 'd0;
    mem[10157] = 'd0;
    mem[10158] = 'd0;
    mem[10159] = 'd856;
    mem[10160] = 'd0;
    mem[10161] = 'd1020;
    mem[10162] = 'd0;
    mem[10163] = 'd0;
    mem[10164] = 'd0;
    mem[10165] = 'd864;
    mem[10166] = 'd0;
    mem[10167] = 'd1020;
    mem[10168] = 'd0;
    mem[10169] = 'd0;
    mem[10170] = 'd0;
    mem[10171] = 'd864;
    mem[10172] = 'd0;
    mem[10173] = 'd1020;
    mem[10174] = 'd0;
    mem[10175] = 'd0;
    mem[10176] = 'd0;
    mem[10177] = 'd864;
    mem[10178] = 'd0;
    mem[10179] = 'd1020;
    mem[10180] = 'd0;
    mem[10181] = 'd0;
    mem[10182] = 'd0;
    mem[10183] = 'd864;
    mem[10184] = 'd0;
    mem[10185] = 'd1020;
    mem[10186] = 'd0;
    mem[10187] = 'd0;
    mem[10188] = 'd0;
    mem[10189] = 'd856;
    mem[10190] = 'd0;
    mem[10191] = 'd1016;
    mem[10192] = 'd0;
    mem[10193] = 'd0;
    mem[10194] = 'd0;
    mem[10195] = 'd812;
    mem[10196] = 'd0;
    mem[10197] = 'd996;
    mem[10198] = 'd0;
    mem[10199] = 'd0;
    mem[10200] = 'd0;
    mem[10201] = 'd572;
    mem[10202] = 'd0;
    mem[10203] = 'd736;
    mem[10204] = 'd0;
    mem[10205] = 'd0;
    mem[10206] = 'd0;
    mem[10207] = 'd292;
    mem[10208] = 'd0;
    mem[10209] = 'd376;
    mem[10210] = 'd0;
    mem[10211] = 'd0;
    mem[10212] = 'd0;
    mem[10213] = 'd188;
    mem[10214] = 'd0;
    mem[10215] = 'd244;
    mem[10216] = 'd0;
    mem[10217] = 'd0;
    mem[10218] = 'd0;
    mem[10219] = 'd148;
    mem[10220] = 'd0;
    mem[10221] = 'd188;
    mem[10222] = 'd0;
    mem[10223] = 'd0;
    mem[10224] = 'd0;
    mem[10225] = 'd176;
    mem[10226] = 'd0;
    mem[10227] = 'd232;
    mem[10228] = 'd0;
    mem[10229] = 'd0;
    mem[10230] = 'd0;
    mem[10231] = 'd276;
    mem[10232] = 'd0;
    mem[10233] = 'd384;
    mem[10234] = 'd0;
    mem[10235] = 'd0;
    mem[10236] = 'd0;
    mem[10237] = 'd428;
    mem[10238] = 'd0;
    mem[10239] = 'd604;
    mem[10240] = 'd0;
    mem[10241] = 'd0;
    mem[10242] = 'd0;
    mem[10243] = 'd632;
    mem[10244] = 'd0;
    mem[10245] = 'd900;
    mem[10246] = 'd0;
    mem[10247] = 'd0;
    mem[10248] = 'd0;
    mem[10249] = 'd692;
    mem[10250] = 'd0;
    mem[10251] = 'd956;
    mem[10252] = 'd0;
    mem[10253] = 'd0;
    mem[10254] = 'd0;
    mem[10255] = 'd724;
    mem[10256] = 'd0;
    mem[10257] = 'd1004;
    mem[10258] = 'd0;
    mem[10259] = 'd0;
    mem[10260] = 'd0;
    mem[10261] = 'd700;
    mem[10262] = 'd0;
    mem[10263] = 'd1004;
    mem[10264] = 'd0;
    mem[10265] = 'd0;
    mem[10266] = 'd0;
    mem[10267] = 'd636;
    mem[10268] = 'd0;
    mem[10269] = 'd964;
    mem[10270] = 'd0;
    mem[10271] = 'd0;
    mem[10272] = 'd0;
    mem[10273] = 'd548;
    mem[10274] = 'd0;
    mem[10275] = 'd912;
    mem[10276] = 'd0;
    mem[10277] = 'd0;
    mem[10278] = 'd0;
    mem[10279] = 'd568;
    mem[10280] = 'd0;
    mem[10281] = 'd872;
    mem[10282] = 'd0;
    mem[10283] = 'd0;
    mem[10284] = 'd0;
    mem[10285] = 'd1020;
    mem[10286] = 'd0;
    mem[10287] = 'd1020;
    mem[10288] = 'd0;
    mem[10289] = 'd0;
    mem[10290] = 'd0;
    mem[10291] = 'd1020;
    mem[10292] = 'd0;
    mem[10293] = 'd1020;
    mem[10294] = 'd0;
    mem[10295] = 'd0;
    mem[10296] = 'd0;
    mem[10297] = 'd0;
    mem[10298] = 'd1020;
    mem[10299] = 'd0;
    mem[10300] = 'd1020;
    mem[10301] = 'd0;
    mem[10302] = 'd0;
    mem[10303] = 'd0;
    mem[10304] = 'd448;
    mem[10305] = 'd0;
    mem[10306] = 'd676;
    mem[10307] = 'd0;
    mem[10308] = 'd0;
    mem[10309] = 'd0;
    mem[10310] = 'd20;
    mem[10311] = 'd0;
    mem[10312] = 'd516;
    mem[10313] = 'd0;
    mem[10314] = 'd0;
    mem[10315] = 'd0;
    mem[10316] = 'd44;
    mem[10317] = 'd0;
    mem[10318] = 'd612;
    mem[10319] = 'd0;
    mem[10320] = 'd0;
    mem[10321] = 'd0;
    mem[10322] = 'd68;
    mem[10323] = 'd0;
    mem[10324] = 'd684;
    mem[10325] = 'd0;
    mem[10326] = 'd0;
    mem[10327] = 'd0;
    mem[10328] = 'd120;
    mem[10329] = 'd0;
    mem[10330] = 'd720;
    mem[10331] = 'd0;
    mem[10332] = 'd0;
    mem[10333] = 'd0;
    mem[10334] = 'd172;
    mem[10335] = 'd0;
    mem[10336] = 'd744;
    mem[10337] = 'd0;
    mem[10338] = 'd0;
    mem[10339] = 'd0;
    mem[10340] = 'd188;
    mem[10341] = 'd0;
    mem[10342] = 'd760;
    mem[10343] = 'd0;
    mem[10344] = 'd0;
    mem[10345] = 'd0;
    mem[10346] = 'd180;
    mem[10347] = 'd0;
    mem[10348] = 'd760;
    mem[10349] = 'd0;
    mem[10350] = 'd0;
    mem[10351] = 'd0;
    mem[10352] = 'd172;
    mem[10353] = 'd0;
    mem[10354] = 'd756;
    mem[10355] = 'd0;
    mem[10356] = 'd0;
    mem[10357] = 'd0;
    mem[10358] = 'd160;
    mem[10359] = 'd0;
    mem[10360] = 'd756;
    mem[10361] = 'd0;
    mem[10362] = 'd0;
    mem[10363] = 'd0;
    mem[10364] = 'd164;
    mem[10365] = 'd0;
    mem[10366] = 'd768;
    mem[10367] = 'd0;
    mem[10368] = 'd0;
    mem[10369] = 'd0;
    mem[10370] = 'd176;
    mem[10371] = 'd0;
    mem[10372] = 'd788;
    mem[10373] = 'd0;
    mem[10374] = 'd0;
    mem[10375] = 'd0;
    mem[10376] = 'd196;
    mem[10377] = 'd0;
    mem[10378] = 'd812;
    mem[10379] = 'd0;
    mem[10380] = 'd0;
    mem[10381] = 'd0;
    mem[10382] = 'd204;
    mem[10383] = 'd0;
    mem[10384] = 'd836;
    mem[10385] = 'd0;
    mem[10386] = 'd0;
    mem[10387] = 'd0;
    mem[10388] = 'd208;
    mem[10389] = 'd0;
    mem[10390] = 'd844;
    mem[10391] = 'd0;
    mem[10392] = 'd0;
    mem[10393] = 'd0;
    mem[10394] = 'd212;
    mem[10395] = 'd0;
    mem[10396] = 'd848;
    mem[10397] = 'd0;
    mem[10398] = 'd0;
    mem[10399] = 'd0;
    mem[10400] = 'd208;
    mem[10401] = 'd0;
    mem[10402] = 'd852;
    mem[10403] = 'd0;
    mem[10404] = 'd0;
    mem[10405] = 'd0;
    mem[10406] = 'd208;
    mem[10407] = 'd0;
    mem[10408] = 'd852;
    mem[10409] = 'd0;
    mem[10410] = 'd0;
    mem[10411] = 'd0;
    mem[10412] = 'd208;
    mem[10413] = 'd0;
    mem[10414] = 'd852;
    mem[10415] = 'd0;
    mem[10416] = 'd0;
    mem[10417] = 'd0;
    mem[10418] = 'd208;
    mem[10419] = 'd0;
    mem[10420] = 'd852;
    mem[10421] = 'd0;
    mem[10422] = 'd0;
    mem[10423] = 'd0;
    mem[10424] = 'd208;
    mem[10425] = 'd0;
    mem[10426] = 'd852;
    mem[10427] = 'd0;
    mem[10428] = 'd0;
    mem[10429] = 'd0;
    mem[10430] = 'd208;
    mem[10431] = 'd0;
    mem[10432] = 'd844;
    mem[10433] = 'd0;
    mem[10434] = 'd0;
    mem[10435] = 'd0;
    mem[10436] = 'd200;
    mem[10437] = 'd0;
    mem[10438] = 'd832;
    mem[10439] = 'd0;
    mem[10440] = 'd0;
    mem[10441] = 'd0;
    mem[10442] = 'd184;
    mem[10443] = 'd0;
    mem[10444] = 'd800;
    mem[10445] = 'd0;
    mem[10446] = 'd0;
    mem[10447] = 'd0;
    mem[10448] = 'd160;
    mem[10449] = 'd0;
    mem[10450] = 'd764;
    mem[10451] = 'd0;
    mem[10452] = 'd0;
    mem[10453] = 'd0;
    mem[10454] = 'd148;
    mem[10455] = 'd0;
    mem[10456] = 'd744;
    mem[10457] = 'd0;
    mem[10458] = 'd0;
    mem[10459] = 'd0;
    mem[10460] = 'd148;
    mem[10461] = 'd0;
    mem[10462] = 'd736;
    mem[10463] = 'd0;
    mem[10464] = 'd0;
    mem[10465] = 'd0;
    mem[10466] = 'd160;
    mem[10467] = 'd0;
    mem[10468] = 'd740;
    mem[10469] = 'd0;
    mem[10470] = 'd0;
    mem[10471] = 'd0;
    mem[10472] = 'd172;
    mem[10473] = 'd0;
    mem[10474] = 'd748;
    mem[10475] = 'd0;
    mem[10476] = 'd0;
    mem[10477] = 'd0;
    mem[10478] = 'd188;
    mem[10479] = 'd0;
    mem[10480] = 'd756;
    mem[10481] = 'd0;
    mem[10482] = 'd0;
    mem[10483] = 'd0;
    mem[10484] = 'd172;
    mem[10485] = 'd0;
    mem[10486] = 'd748;
    mem[10487] = 'd0;
    mem[10488] = 'd0;
    mem[10489] = 'd0;
    mem[10490] = 'd120;
    mem[10491] = 'd0;
    mem[10492] = 'd724;
    mem[10493] = 'd0;
    mem[10494] = 'd0;
    mem[10495] = 'd0;
    mem[10496] = 'd72;
    mem[10497] = 'd0;
    mem[10498] = 'd684;
    mem[10499] = 'd0;
    mem[10500] = 'd0;
    mem[10501] = 'd0;
    mem[10502] = 'd48;
    mem[10503] = 'd0;
    mem[10504] = 'd616;
    mem[10505] = 'd0;
    mem[10506] = 'd0;
    mem[10507] = 'd0;
    mem[10508] = 'd24;
    mem[10509] = 'd0;
    mem[10510] = 'd524;
    mem[10511] = 'd0;
    mem[10512] = 'd0;
    mem[10513] = 'd0;
    mem[10514] = 'd404;
    mem[10515] = 'd0;
    mem[10516] = 'd660;
    mem[10517] = 'd0;
    mem[10518] = 'd0;
    mem[10519] = 'd0;
    mem[10520] = 'd1020;
    mem[10521] = 'd0;
    mem[10522] = 'd1020;
    mem[10523] = 'd0;
    mem[10524] = 'd0;
    mem[10525] = 'd0;
    mem[10526] = 'd1020;
    mem[10527] = 'd0;
    mem[10528] = 'd1020;
    mem[10529] = 'd0;
    mem[10530] = 'd0;
    mem[10531] = 'd1020;
    mem[10532] = 'd0;
    mem[10533] = 'd1020;
    mem[10534] = 'd0;
    mem[10535] = 'd0;
    mem[10536] = 'd0;
    mem[10537] = 'd676;
    mem[10538] = 'd0;
    mem[10539] = 'd900;
    mem[10540] = 'd0;
    mem[10541] = 'd0;
    mem[10542] = 'd0;
    mem[10543] = 'd516;
    mem[10544] = 'd0;
    mem[10545] = 'd884;
    mem[10546] = 'd0;
    mem[10547] = 'd0;
    mem[10548] = 'd0;
    mem[10549] = 'd612;
    mem[10550] = 'd0;
    mem[10551] = 'd944;
    mem[10552] = 'd0;
    mem[10553] = 'd0;
    mem[10554] = 'd0;
    mem[10555] = 'd684;
    mem[10556] = 'd0;
    mem[10557] = 'd996;
    mem[10558] = 'd0;
    mem[10559] = 'd0;
    mem[10560] = 'd0;
    mem[10561] = 'd720;
    mem[10562] = 'd0;
    mem[10563] = 'd1012;
    mem[10564] = 'd0;
    mem[10565] = 'd0;
    mem[10566] = 'd0;
    mem[10567] = 'd744;
    mem[10568] = 'd0;
    mem[10569] = 'd1016;
    mem[10570] = 'd0;
    mem[10571] = 'd0;
    mem[10572] = 'd0;
    mem[10573] = 'd760;
    mem[10574] = 'd0;
    mem[10575] = 'd1012;
    mem[10576] = 'd0;
    mem[10577] = 'd0;
    mem[10578] = 'd0;
    mem[10579] = 'd760;
    mem[10580] = 'd0;
    mem[10581] = 'd1000;
    mem[10582] = 'd0;
    mem[10583] = 'd0;
    mem[10584] = 'd0;
    mem[10585] = 'd756;
    mem[10586] = 'd0;
    mem[10587] = 'd988;
    mem[10588] = 'd0;
    mem[10589] = 'd0;
    mem[10590] = 'd0;
    mem[10591] = 'd756;
    mem[10592] = 'd0;
    mem[10593] = 'd988;
    mem[10594] = 'd0;
    mem[10595] = 'd0;
    mem[10596] = 'd0;
    mem[10597] = 'd768;
    mem[10598] = 'd0;
    mem[10599] = 'd992;
    mem[10600] = 'd0;
    mem[10601] = 'd0;
    mem[10602] = 'd0;
    mem[10603] = 'd788;
    mem[10604] = 'd0;
    mem[10605] = 'd1000;
    mem[10606] = 'd0;
    mem[10607] = 'd0;
    mem[10608] = 'd0;
    mem[10609] = 'd812;
    mem[10610] = 'd0;
    mem[10611] = 'd1008;
    mem[10612] = 'd0;
    mem[10613] = 'd0;
    mem[10614] = 'd0;
    mem[10615] = 'd836;
    mem[10616] = 'd0;
    mem[10617] = 'd1016;
    mem[10618] = 'd0;
    mem[10619] = 'd0;
    mem[10620] = 'd0;
    mem[10621] = 'd844;
    mem[10622] = 'd0;
    mem[10623] = 'd1020;
    mem[10624] = 'd0;
    mem[10625] = 'd0;
    mem[10626] = 'd0;
    mem[10627] = 'd848;
    mem[10628] = 'd0;
    mem[10629] = 'd1020;
    mem[10630] = 'd0;
    mem[10631] = 'd0;
    mem[10632] = 'd0;
    mem[10633] = 'd852;
    mem[10634] = 'd0;
    mem[10635] = 'd1020;
    mem[10636] = 'd0;
    mem[10637] = 'd0;
    mem[10638] = 'd0;
    mem[10639] = 'd852;
    mem[10640] = 'd0;
    mem[10641] = 'd1020;
    mem[10642] = 'd0;
    mem[10643] = 'd0;
    mem[10644] = 'd0;
    mem[10645] = 'd852;
    mem[10646] = 'd0;
    mem[10647] = 'd1020;
    mem[10648] = 'd0;
    mem[10649] = 'd0;
    mem[10650] = 'd0;
    mem[10651] = 'd852;
    mem[10652] = 'd0;
    mem[10653] = 'd1020;
    mem[10654] = 'd0;
    mem[10655] = 'd0;
    mem[10656] = 'd0;
    mem[10657] = 'd852;
    mem[10658] = 'd0;
    mem[10659] = 'd1020;
    mem[10660] = 'd0;
    mem[10661] = 'd0;
    mem[10662] = 'd0;
    mem[10663] = 'd844;
    mem[10664] = 'd0;
    mem[10665] = 'd1020;
    mem[10666] = 'd0;
    mem[10667] = 'd0;
    mem[10668] = 'd0;
    mem[10669] = 'd832;
    mem[10670] = 'd0;
    mem[10671] = 'd1012;
    mem[10672] = 'd0;
    mem[10673] = 'd0;
    mem[10674] = 'd0;
    mem[10675] = 'd800;
    mem[10676] = 'd0;
    mem[10677] = 'd996;
    mem[10678] = 'd0;
    mem[10679] = 'd0;
    mem[10680] = 'd0;
    mem[10681] = 'd764;
    mem[10682] = 'd0;
    mem[10683] = 'd984;
    mem[10684] = 'd0;
    mem[10685] = 'd0;
    mem[10686] = 'd0;
    mem[10687] = 'd744;
    mem[10688] = 'd0;
    mem[10689] = 'd976;
    mem[10690] = 'd0;
    mem[10691] = 'd0;
    mem[10692] = 'd0;
    mem[10693] = 'd736;
    mem[10694] = 'd0;
    mem[10695] = 'd972;
    mem[10696] = 'd0;
    mem[10697] = 'd0;
    mem[10698] = 'd0;
    mem[10699] = 'd740;
    mem[10700] = 'd0;
    mem[10701] = 'd976;
    mem[10702] = 'd0;
    mem[10703] = 'd0;
    mem[10704] = 'd0;
    mem[10705] = 'd748;
    mem[10706] = 'd0;
    mem[10707] = 'd992;
    mem[10708] = 'd0;
    mem[10709] = 'd0;
    mem[10710] = 'd0;
    mem[10711] = 'd756;
    mem[10712] = 'd0;
    mem[10713] = 'd1008;
    mem[10714] = 'd0;
    mem[10715] = 'd0;
    mem[10716] = 'd0;
    mem[10717] = 'd748;
    mem[10718] = 'd0;
    mem[10719] = 'd1016;
    mem[10720] = 'd0;
    mem[10721] = 'd0;
    mem[10722] = 'd0;
    mem[10723] = 'd724;
    mem[10724] = 'd0;
    mem[10725] = 'd1012;
    mem[10726] = 'd0;
    mem[10727] = 'd0;
    mem[10728] = 'd0;
    mem[10729] = 'd684;
    mem[10730] = 'd0;
    mem[10731] = 'd996;
    mem[10732] = 'd0;
    mem[10733] = 'd0;
    mem[10734] = 'd0;
    mem[10735] = 'd616;
    mem[10736] = 'd0;
    mem[10737] = 'd948;
    mem[10738] = 'd0;
    mem[10739] = 'd0;
    mem[10740] = 'd0;
    mem[10741] = 'd524;
    mem[10742] = 'd0;
    mem[10743] = 'd892;
    mem[10744] = 'd0;
    mem[10745] = 'd0;
    mem[10746] = 'd0;
    mem[10747] = 'd660;
    mem[10748] = 'd0;
    mem[10749] = 'd892;
    mem[10750] = 'd0;
    mem[10751] = 'd0;
    mem[10752] = 'd0;
    mem[10753] = 'd1020;
    mem[10754] = 'd0;
    mem[10755] = 'd1020;
    mem[10756] = 'd0;
    mem[10757] = 'd0;
    mem[10758] = 'd0;
    mem[10759] = 'd1020;
    mem[10760] = 'd0;
    mem[10761] = 'd1020;
    mem[10762] = 'd0;
    mem[10763] = 'd0;
    mem[10764] = 'd0;
    mem[10765] = 'd0;
    mem[10766] = 'd1020;
    mem[10767] = 'd0;
    mem[10768] = 'd1020;
    mem[10769] = 'd0;
    mem[10770] = 'd0;
    mem[10771] = 'd0;
    mem[10772] = 'd676;
    mem[10773] = 'd0;
    mem[10774] = 'd808;
    mem[10775] = 'd0;
    mem[10776] = 'd0;
    mem[10777] = 'd0;
    mem[10778] = 'd16;
    mem[10779] = 'd0;
    mem[10780] = 'd488;
    mem[10781] = 'd0;
    mem[10782] = 'd0;
    mem[10783] = 'd0;
    mem[10784] = 'd40;
    mem[10785] = 'd0;
    mem[10786] = 'd584;
    mem[10787] = 'd0;
    mem[10788] = 'd0;
    mem[10789] = 'd0;
    mem[10790] = 'd64;
    mem[10791] = 'd0;
    mem[10792] = 'd660;
    mem[10793] = 'd0;
    mem[10794] = 'd0;
    mem[10795] = 'd0;
    mem[10796] = 'd92;
    mem[10797] = 'd0;
    mem[10798] = 'd704;
    mem[10799] = 'd0;
    mem[10800] = 'd0;
    mem[10801] = 'd0;
    mem[10802] = 'd140;
    mem[10803] = 'd0;
    mem[10804] = 'd732;
    mem[10805] = 'd0;
    mem[10806] = 'd0;
    mem[10807] = 'd0;
    mem[10808] = 'd184;
    mem[10809] = 'd0;
    mem[10810] = 'd756;
    mem[10811] = 'd0;
    mem[10812] = 'd0;
    mem[10813] = 'd0;
    mem[10814] = 'd208;
    mem[10815] = 'd0;
    mem[10816] = 'd772;
    mem[10817] = 'd0;
    mem[10818] = 'd0;
    mem[10819] = 'd0;
    mem[10820] = 'd212;
    mem[10821] = 'd0;
    mem[10822] = 'd784;
    mem[10823] = 'd0;
    mem[10824] = 'd0;
    mem[10825] = 'd0;
    mem[10826] = 'd200;
    mem[10827] = 'd0;
    mem[10828] = 'd780;
    mem[10829] = 'd0;
    mem[10830] = 'd0;
    mem[10831] = 'd0;
    mem[10832] = 'd204;
    mem[10833] = 'd0;
    mem[10834] = 'd800;
    mem[10835] = 'd0;
    mem[10836] = 'd0;
    mem[10837] = 'd0;
    mem[10838] = 'd212;
    mem[10839] = 'd0;
    mem[10840] = 'd816;
    mem[10841] = 'd0;
    mem[10842] = 'd0;
    mem[10843] = 'd0;
    mem[10844] = 'd216;
    mem[10845] = 'd0;
    mem[10846] = 'd824;
    mem[10847] = 'd0;
    mem[10848] = 'd0;
    mem[10849] = 'd0;
    mem[10850] = 'd216;
    mem[10851] = 'd0;
    mem[10852] = 'd832;
    mem[10853] = 'd0;
    mem[10854] = 'd0;
    mem[10855] = 'd0;
    mem[10856] = 'd216;
    mem[10857] = 'd0;
    mem[10858] = 'd836;
    mem[10859] = 'd0;
    mem[10860] = 'd0;
    mem[10861] = 'd0;
    mem[10862] = 'd216;
    mem[10863] = 'd0;
    mem[10864] = 'd836;
    mem[10865] = 'd0;
    mem[10866] = 'd0;
    mem[10867] = 'd0;
    mem[10868] = 'd216;
    mem[10869] = 'd0;
    mem[10870] = 'd840;
    mem[10871] = 'd0;
    mem[10872] = 'd0;
    mem[10873] = 'd0;
    mem[10874] = 'd220;
    mem[10875] = 'd0;
    mem[10876] = 'd840;
    mem[10877] = 'd0;
    mem[10878] = 'd0;
    mem[10879] = 'd0;
    mem[10880] = 'd216;
    mem[10881] = 'd0;
    mem[10882] = 'd844;
    mem[10883] = 'd0;
    mem[10884] = 'd0;
    mem[10885] = 'd0;
    mem[10886] = 'd216;
    mem[10887] = 'd0;
    mem[10888] = 'd840;
    mem[10889] = 'd0;
    mem[10890] = 'd0;
    mem[10891] = 'd0;
    mem[10892] = 'd216;
    mem[10893] = 'd0;
    mem[10894] = 'd836;
    mem[10895] = 'd0;
    mem[10896] = 'd0;
    mem[10897] = 'd0;
    mem[10898] = 'd216;
    mem[10899] = 'd0;
    mem[10900] = 'd836;
    mem[10901] = 'd0;
    mem[10902] = 'd0;
    mem[10903] = 'd0;
    mem[10904] = 'd216;
    mem[10905] = 'd0;
    mem[10906] = 'd832;
    mem[10907] = 'd0;
    mem[10908] = 'd0;
    mem[10909] = 'd0;
    mem[10910] = 'd216;
    mem[10911] = 'd0;
    mem[10912] = 'd824;
    mem[10913] = 'd0;
    mem[10914] = 'd0;
    mem[10915] = 'd0;
    mem[10916] = 'd216;
    mem[10917] = 'd0;
    mem[10918] = 'd820;
    mem[10919] = 'd0;
    mem[10920] = 'd0;
    mem[10921] = 'd0;
    mem[10922] = 'd208;
    mem[10923] = 'd0;
    mem[10924] = 'd800;
    mem[10925] = 'd0;
    mem[10926] = 'd0;
    mem[10927] = 'd0;
    mem[10928] = 'd200;
    mem[10929] = 'd0;
    mem[10930] = 'd776;
    mem[10931] = 'd0;
    mem[10932] = 'd0;
    mem[10933] = 'd0;
    mem[10934] = 'd212;
    mem[10935] = 'd0;
    mem[10936] = 'd784;
    mem[10937] = 'd0;
    mem[10938] = 'd0;
    mem[10939] = 'd0;
    mem[10940] = 'd208;
    mem[10941] = 'd0;
    mem[10942] = 'd772;
    mem[10943] = 'd0;
    mem[10944] = 'd0;
    mem[10945] = 'd0;
    mem[10946] = 'd184;
    mem[10947] = 'd0;
    mem[10948] = 'd756;
    mem[10949] = 'd0;
    mem[10950] = 'd0;
    mem[10951] = 'd0;
    mem[10952] = 'd144;
    mem[10953] = 'd0;
    mem[10954] = 'd732;
    mem[10955] = 'd0;
    mem[10956] = 'd0;
    mem[10957] = 'd0;
    mem[10958] = 'd92;
    mem[10959] = 'd0;
    mem[10960] = 'd708;
    mem[10961] = 'd0;
    mem[10962] = 'd0;
    mem[10963] = 'd0;
    mem[10964] = 'd64;
    mem[10965] = 'd0;
    mem[10966] = 'd660;
    mem[10967] = 'd0;
    mem[10968] = 'd0;
    mem[10969] = 'd0;
    mem[10970] = 'd44;
    mem[10971] = 'd0;
    mem[10972] = 'd588;
    mem[10973] = 'd0;
    mem[10974] = 'd0;
    mem[10975] = 'd0;
    mem[10976] = 'd16;
    mem[10977] = 'd0;
    mem[10978] = 'd492;
    mem[10979] = 'd0;
    mem[10980] = 'd0;
    mem[10981] = 'd0;
    mem[10982] = 'd636;
    mem[10983] = 'd0;
    mem[10984] = 'd788;
    mem[10985] = 'd0;
    mem[10986] = 'd0;
    mem[10987] = 'd0;
    mem[10988] = 'd1020;
    mem[10989] = 'd0;
    mem[10990] = 'd1020;
    mem[10991] = 'd0;
    mem[10992] = 'd0;
    mem[10993] = 'd0;
    mem[10994] = 'd1020;
    mem[10995] = 'd0;
    mem[10996] = 'd1020;
    mem[10997] = 'd0;
    mem[10998] = 'd0;
    mem[10999] = 'd1020;
    mem[11000] = 'd0;
    mem[11001] = 'd1020;
    mem[11002] = 'd0;
    mem[11003] = 'd0;
    mem[11004] = 'd0;
    mem[11005] = 'd808;
    mem[11006] = 'd0;
    mem[11007] = 'd936;
    mem[11008] = 'd0;
    mem[11009] = 'd0;
    mem[11010] = 'd0;
    mem[11011] = 'd488;
    mem[11012] = 'd0;
    mem[11013] = 'd860;
    mem[11014] = 'd0;
    mem[11015] = 'd0;
    mem[11016] = 'd0;
    mem[11017] = 'd584;
    mem[11018] = 'd0;
    mem[11019] = 'd924;
    mem[11020] = 'd0;
    mem[11021] = 'd0;
    mem[11022] = 'd0;
    mem[11023] = 'd660;
    mem[11024] = 'd0;
    mem[11025] = 'd976;
    mem[11026] = 'd0;
    mem[11027] = 'd0;
    mem[11028] = 'd0;
    mem[11029] = 'd704;
    mem[11030] = 'd0;
    mem[11031] = 'd1008;
    mem[11032] = 'd0;
    mem[11033] = 'd0;
    mem[11034] = 'd0;
    mem[11035] = 'd732;
    mem[11036] = 'd0;
    mem[11037] = 'd1016;
    mem[11038] = 'd0;
    mem[11039] = 'd0;
    mem[11040] = 'd0;
    mem[11041] = 'd756;
    mem[11042] = 'd0;
    mem[11043] = 'd1020;
    mem[11044] = 'd0;
    mem[11045] = 'd0;
    mem[11046] = 'd0;
    mem[11047] = 'd772;
    mem[11048] = 'd0;
    mem[11049] = 'd1020;
    mem[11050] = 'd0;
    mem[11051] = 'd0;
    mem[11052] = 'd0;
    mem[11053] = 'd784;
    mem[11054] = 'd0;
    mem[11055] = 'd1020;
    mem[11056] = 'd0;
    mem[11057] = 'd0;
    mem[11058] = 'd0;
    mem[11059] = 'd780;
    mem[11060] = 'd0;
    mem[11061] = 'd1008;
    mem[11062] = 'd0;
    mem[11063] = 'd0;
    mem[11064] = 'd0;
    mem[11065] = 'd800;
    mem[11066] = 'd0;
    mem[11067] = 'd1012;
    mem[11068] = 'd0;
    mem[11069] = 'd0;
    mem[11070] = 'd0;
    mem[11071] = 'd816;
    mem[11072] = 'd0;
    mem[11073] = 'd1020;
    mem[11074] = 'd0;
    mem[11075] = 'd0;
    mem[11076] = 'd0;
    mem[11077] = 'd824;
    mem[11078] = 'd0;
    mem[11079] = 'd1020;
    mem[11080] = 'd0;
    mem[11081] = 'd0;
    mem[11082] = 'd0;
    mem[11083] = 'd832;
    mem[11084] = 'd0;
    mem[11085] = 'd1020;
    mem[11086] = 'd0;
    mem[11087] = 'd0;
    mem[11088] = 'd0;
    mem[11089] = 'd836;
    mem[11090] = 'd0;
    mem[11091] = 'd1020;
    mem[11092] = 'd0;
    mem[11093] = 'd0;
    mem[11094] = 'd0;
    mem[11095] = 'd836;
    mem[11096] = 'd0;
    mem[11097] = 'd1020;
    mem[11098] = 'd0;
    mem[11099] = 'd0;
    mem[11100] = 'd0;
    mem[11101] = 'd840;
    mem[11102] = 'd0;
    mem[11103] = 'd1020;
    mem[11104] = 'd0;
    mem[11105] = 'd0;
    mem[11106] = 'd0;
    mem[11107] = 'd840;
    mem[11108] = 'd0;
    mem[11109] = 'd1020;
    mem[11110] = 'd0;
    mem[11111] = 'd0;
    mem[11112] = 'd0;
    mem[11113] = 'd844;
    mem[11114] = 'd0;
    mem[11115] = 'd1020;
    mem[11116] = 'd0;
    mem[11117] = 'd0;
    mem[11118] = 'd0;
    mem[11119] = 'd840;
    mem[11120] = 'd0;
    mem[11121] = 'd1020;
    mem[11122] = 'd0;
    mem[11123] = 'd0;
    mem[11124] = 'd0;
    mem[11125] = 'd836;
    mem[11126] = 'd0;
    mem[11127] = 'd1020;
    mem[11128] = 'd0;
    mem[11129] = 'd0;
    mem[11130] = 'd0;
    mem[11131] = 'd836;
    mem[11132] = 'd0;
    mem[11133] = 'd1020;
    mem[11134] = 'd0;
    mem[11135] = 'd0;
    mem[11136] = 'd0;
    mem[11137] = 'd832;
    mem[11138] = 'd0;
    mem[11139] = 'd1020;
    mem[11140] = 'd0;
    mem[11141] = 'd0;
    mem[11142] = 'd0;
    mem[11143] = 'd824;
    mem[11144] = 'd0;
    mem[11145] = 'd1020;
    mem[11146] = 'd0;
    mem[11147] = 'd0;
    mem[11148] = 'd0;
    mem[11149] = 'd820;
    mem[11150] = 'd0;
    mem[11151] = 'd1020;
    mem[11152] = 'd0;
    mem[11153] = 'd0;
    mem[11154] = 'd0;
    mem[11155] = 'd800;
    mem[11156] = 'd0;
    mem[11157] = 'd1016;
    mem[11158] = 'd0;
    mem[11159] = 'd0;
    mem[11160] = 'd0;
    mem[11161] = 'd776;
    mem[11162] = 'd0;
    mem[11163] = 'd1012;
    mem[11164] = 'd0;
    mem[11165] = 'd0;
    mem[11166] = 'd0;
    mem[11167] = 'd784;
    mem[11168] = 'd0;
    mem[11169] = 'd1020;
    mem[11170] = 'd0;
    mem[11171] = 'd0;
    mem[11172] = 'd0;
    mem[11173] = 'd772;
    mem[11174] = 'd0;
    mem[11175] = 'd1020;
    mem[11176] = 'd0;
    mem[11177] = 'd0;
    mem[11178] = 'd0;
    mem[11179] = 'd756;
    mem[11180] = 'd0;
    mem[11181] = 'd1020;
    mem[11182] = 'd0;
    mem[11183] = 'd0;
    mem[11184] = 'd0;
    mem[11185] = 'd732;
    mem[11186] = 'd0;
    mem[11187] = 'd1016;
    mem[11188] = 'd0;
    mem[11189] = 'd0;
    mem[11190] = 'd0;
    mem[11191] = 'd708;
    mem[11192] = 'd0;
    mem[11193] = 'd1008;
    mem[11194] = 'd0;
    mem[11195] = 'd0;
    mem[11196] = 'd0;
    mem[11197] = 'd660;
    mem[11198] = 'd0;
    mem[11199] = 'd976;
    mem[11200] = 'd0;
    mem[11201] = 'd0;
    mem[11202] = 'd0;
    mem[11203] = 'd588;
    mem[11204] = 'd0;
    mem[11205] = 'd928;
    mem[11206] = 'd0;
    mem[11207] = 'd0;
    mem[11208] = 'd0;
    mem[11209] = 'd492;
    mem[11210] = 'd0;
    mem[11211] = 'd864;
    mem[11212] = 'd0;
    mem[11213] = 'd0;
    mem[11214] = 'd0;
    mem[11215] = 'd788;
    mem[11216] = 'd0;
    mem[11217] = 'd928;
    mem[11218] = 'd0;
    mem[11219] = 'd0;
    mem[11220] = 'd0;
    mem[11221] = 'd1020;
    mem[11222] = 'd0;
    mem[11223] = 'd1020;
    mem[11224] = 'd0;
    mem[11225] = 'd0;
    mem[11226] = 'd0;
    mem[11227] = 'd1020;
    mem[11228] = 'd0;
    mem[11229] = 'd1020;
    mem[11230] = 'd0;
    mem[11231] = 'd0;
    mem[11232] = 'd0;
    mem[11233] = 'd0;
    mem[11234] = 'd1020;
    mem[11235] = 'd0;
    mem[11236] = 'd1020;
    mem[11237] = 'd0;
    mem[11238] = 'd0;
    mem[11239] = 'd0;
    mem[11240] = 'd944;
    mem[11241] = 'd0;
    mem[11242] = 'd968;
    mem[11243] = 'd0;
    mem[11244] = 'd0;
    mem[11245] = 'd0;
    mem[11246] = 'd36;
    mem[11247] = 'd0;
    mem[11248] = 'd460;
    mem[11249] = 'd0;
    mem[11250] = 'd0;
    mem[11251] = 'd0;
    mem[11252] = 'd36;
    mem[11253] = 'd0;
    mem[11254] = 'd548;
    mem[11255] = 'd0;
    mem[11256] = 'd0;
    mem[11257] = 'd0;
    mem[11258] = 'd56;
    mem[11259] = 'd0;
    mem[11260] = 'd636;
    mem[11261] = 'd0;
    mem[11262] = 'd0;
    mem[11263] = 'd0;
    mem[11264] = 'd76;
    mem[11265] = 'd0;
    mem[11266] = 'd684;
    mem[11267] = 'd0;
    mem[11268] = 'd0;
    mem[11269] = 'd0;
    mem[11270] = 'd108;
    mem[11271] = 'd0;
    mem[11272] = 'd716;
    mem[11273] = 'd0;
    mem[11274] = 'd0;
    mem[11275] = 'd0;
    mem[11276] = 'd156;
    mem[11277] = 'd0;
    mem[11278] = 'd740;
    mem[11279] = 'd0;
    mem[11280] = 'd0;
    mem[11281] = 'd0;
    mem[11282] = 'd196;
    mem[11283] = 'd0;
    mem[11284] = 'd756;
    mem[11285] = 'd0;
    mem[11286] = 'd0;
    mem[11287] = 'd0;
    mem[11288] = 'd216;
    mem[11289] = 'd0;
    mem[11290] = 'd772;
    mem[11291] = 'd0;
    mem[11292] = 'd0;
    mem[11293] = 'd0;
    mem[11294] = 'd112;
    mem[11295] = 'd0;
    mem[11296] = 'd480;
    mem[11297] = 'd0;
    mem[11298] = 'd0;
    mem[11299] = 'd0;
    mem[11300] = 'd104;
    mem[11301] = 'd0;
    mem[11302] = 'd500;
    mem[11303] = 'd0;
    mem[11304] = 'd0;
    mem[11305] = 'd0;
    mem[11306] = 'd200;
    mem[11307] = 'd0;
    mem[11308] = 'd776;
    mem[11309] = 'd0;
    mem[11310] = 'd0;
    mem[11311] = 'd0;
    mem[11312] = 'd216;
    mem[11313] = 'd0;
    mem[11314] = 'd812;
    mem[11315] = 'd0;
    mem[11316] = 'd0;
    mem[11317] = 'd0;
    mem[11318] = 'd224;
    mem[11319] = 'd0;
    mem[11320] = 'd820;
    mem[11321] = 'd0;
    mem[11322] = 'd0;
    mem[11323] = 'd0;
    mem[11324] = 'd220;
    mem[11325] = 'd0;
    mem[11326] = 'd824;
    mem[11327] = 'd0;
    mem[11328] = 'd0;
    mem[11329] = 'd0;
    mem[11330] = 'd224;
    mem[11331] = 'd0;
    mem[11332] = 'd828;
    mem[11333] = 'd0;
    mem[11334] = 'd0;
    mem[11335] = 'd0;
    mem[11336] = 'd220;
    mem[11337] = 'd0;
    mem[11338] = 'd828;
    mem[11339] = 'd0;
    mem[11340] = 'd0;
    mem[11341] = 'd0;
    mem[11342] = 'd220;
    mem[11343] = 'd0;
    mem[11344] = 'd828;
    mem[11345] = 'd0;
    mem[11346] = 'd0;
    mem[11347] = 'd0;
    mem[11348] = 'd220;
    mem[11349] = 'd0;
    mem[11350] = 'd828;
    mem[11351] = 'd0;
    mem[11352] = 'd0;
    mem[11353] = 'd0;
    mem[11354] = 'd220;
    mem[11355] = 'd0;
    mem[11356] = 'd828;
    mem[11357] = 'd0;
    mem[11358] = 'd0;
    mem[11359] = 'd0;
    mem[11360] = 'd220;
    mem[11361] = 'd0;
    mem[11362] = 'd828;
    mem[11363] = 'd0;
    mem[11364] = 'd0;
    mem[11365] = 'd0;
    mem[11366] = 'd220;
    mem[11367] = 'd0;
    mem[11368] = 'd824;
    mem[11369] = 'd0;
    mem[11370] = 'd0;
    mem[11371] = 'd0;
    mem[11372] = 'd220;
    mem[11373] = 'd0;
    mem[11374] = 'd820;
    mem[11375] = 'd0;
    mem[11376] = 'd0;
    mem[11377] = 'd0;
    mem[11378] = 'd220;
    mem[11379] = 'd0;
    mem[11380] = 'd812;
    mem[11381] = 'd0;
    mem[11382] = 'd0;
    mem[11383] = 'd0;
    mem[11384] = 'd200;
    mem[11385] = 'd0;
    mem[11386] = 'd772;
    mem[11387] = 'd0;
    mem[11388] = 'd0;
    mem[11389] = 'd0;
    mem[11390] = 'd84;
    mem[11391] = 'd0;
    mem[11392] = 'd436;
    mem[11393] = 'd0;
    mem[11394] = 'd0;
    mem[11395] = 'd0;
    mem[11396] = 'd136;
    mem[11397] = 'd0;
    mem[11398] = 'd544;
    mem[11399] = 'd0;
    mem[11400] = 'd0;
    mem[11401] = 'd0;
    mem[11402] = 'd216;
    mem[11403] = 'd0;
    mem[11404] = 'd772;
    mem[11405] = 'd0;
    mem[11406] = 'd0;
    mem[11407] = 'd0;
    mem[11408] = 'd196;
    mem[11409] = 'd0;
    mem[11410] = 'd756;
    mem[11411] = 'd0;
    mem[11412] = 'd0;
    mem[11413] = 'd0;
    mem[11414] = 'd156;
    mem[11415] = 'd0;
    mem[11416] = 'd736;
    mem[11417] = 'd0;
    mem[11418] = 'd0;
    mem[11419] = 'd0;
    mem[11420] = 'd112;
    mem[11421] = 'd0;
    mem[11422] = 'd720;
    mem[11423] = 'd0;
    mem[11424] = 'd0;
    mem[11425] = 'd0;
    mem[11426] = 'd76;
    mem[11427] = 'd0;
    mem[11428] = 'd684;
    mem[11429] = 'd0;
    mem[11430] = 'd0;
    mem[11431] = 'd0;
    mem[11432] = 'd60;
    mem[11433] = 'd0;
    mem[11434] = 'd636;
    mem[11435] = 'd0;
    mem[11436] = 'd0;
    mem[11437] = 'd0;
    mem[11438] = 'd36;
    mem[11439] = 'd0;
    mem[11440] = 'd556;
    mem[11441] = 'd0;
    mem[11442] = 'd0;
    mem[11443] = 'd0;
    mem[11444] = 'd24;
    mem[11445] = 'd0;
    mem[11446] = 'd464;
    mem[11447] = 'd0;
    mem[11448] = 'd0;
    mem[11449] = 'd0;
    mem[11450] = 'd916;
    mem[11451] = 'd0;
    mem[11452] = 'd952;
    mem[11453] = 'd0;
    mem[11454] = 'd0;
    mem[11455] = 'd0;
    mem[11456] = 'd1020;
    mem[11457] = 'd0;
    mem[11458] = 'd1020;
    mem[11459] = 'd0;
    mem[11460] = 'd0;
    mem[11461] = 'd0;
    mem[11462] = 'd1020;
    mem[11463] = 'd0;
    mem[11464] = 'd1020;
    mem[11465] = 'd0;
    mem[11466] = 'd0;
    mem[11467] = 'd1020;
    mem[11468] = 'd0;
    mem[11469] = 'd1020;
    mem[11470] = 'd0;
    mem[11471] = 'd0;
    mem[11472] = 'd0;
    mem[11473] = 'd968;
    mem[11474] = 'd0;
    mem[11475] = 'd996;
    mem[11476] = 'd0;
    mem[11477] = 'd0;
    mem[11478] = 'd0;
    mem[11479] = 'd460;
    mem[11480] = 'd0;
    mem[11481] = 'd832;
    mem[11482] = 'd0;
    mem[11483] = 'd0;
    mem[11484] = 'd0;
    mem[11485] = 'd548;
    mem[11486] = 'd0;
    mem[11487] = 'd896;
    mem[11488] = 'd0;
    mem[11489] = 'd0;
    mem[11490] = 'd0;
    mem[11491] = 'd636;
    mem[11492] = 'd0;
    mem[11493] = 'd956;
    mem[11494] = 'd0;
    mem[11495] = 'd0;
    mem[11496] = 'd0;
    mem[11497] = 'd684;
    mem[11498] = 'd0;
    mem[11499] = 'd996;
    mem[11500] = 'd0;
    mem[11501] = 'd0;
    mem[11502] = 'd0;
    mem[11503] = 'd716;
    mem[11504] = 'd0;
    mem[11505] = 'd1012;
    mem[11506] = 'd0;
    mem[11507] = 'd0;
    mem[11508] = 'd0;
    mem[11509] = 'd740;
    mem[11510] = 'd0;
    mem[11511] = 'd1016;
    mem[11512] = 'd0;
    mem[11513] = 'd0;
    mem[11514] = 'd0;
    mem[11515] = 'd756;
    mem[11516] = 'd0;
    mem[11517] = 'd1020;
    mem[11518] = 'd0;
    mem[11519] = 'd0;
    mem[11520] = 'd0;
    mem[11521] = 'd772;
    mem[11522] = 'd0;
    mem[11523] = 'd1020;
    mem[11524] = 'd0;
    mem[11525] = 'd0;
    mem[11526] = 'd0;
    mem[11527] = 'd480;
    mem[11528] = 'd0;
    mem[11529] = 'd704;
    mem[11530] = 'd0;
    mem[11531] = 'd0;
    mem[11532] = 'd0;
    mem[11533] = 'd500;
    mem[11534] = 'd0;
    mem[11535] = 'd748;
    mem[11536] = 'd0;
    mem[11537] = 'd0;
    mem[11538] = 'd0;
    mem[11539] = 'd776;
    mem[11540] = 'd0;
    mem[11541] = 'd1000;
    mem[11542] = 'd0;
    mem[11543] = 'd0;
    mem[11544] = 'd0;
    mem[11545] = 'd812;
    mem[11546] = 'd0;
    mem[11547] = 'd1020;
    mem[11548] = 'd0;
    mem[11549] = 'd0;
    mem[11550] = 'd0;
    mem[11551] = 'd820;
    mem[11552] = 'd0;
    mem[11553] = 'd1020;
    mem[11554] = 'd0;
    mem[11555] = 'd0;
    mem[11556] = 'd0;
    mem[11557] = 'd824;
    mem[11558] = 'd0;
    mem[11559] = 'd1020;
    mem[11560] = 'd0;
    mem[11561] = 'd0;
    mem[11562] = 'd0;
    mem[11563] = 'd828;
    mem[11564] = 'd0;
    mem[11565] = 'd1020;
    mem[11566] = 'd0;
    mem[11567] = 'd0;
    mem[11568] = 'd0;
    mem[11569] = 'd828;
    mem[11570] = 'd0;
    mem[11571] = 'd1020;
    mem[11572] = 'd0;
    mem[11573] = 'd0;
    mem[11574] = 'd0;
    mem[11575] = 'd828;
    mem[11576] = 'd0;
    mem[11577] = 'd1020;
    mem[11578] = 'd0;
    mem[11579] = 'd0;
    mem[11580] = 'd0;
    mem[11581] = 'd828;
    mem[11582] = 'd0;
    mem[11583] = 'd1020;
    mem[11584] = 'd0;
    mem[11585] = 'd0;
    mem[11586] = 'd0;
    mem[11587] = 'd828;
    mem[11588] = 'd0;
    mem[11589] = 'd1020;
    mem[11590] = 'd0;
    mem[11591] = 'd0;
    mem[11592] = 'd0;
    mem[11593] = 'd828;
    mem[11594] = 'd0;
    mem[11595] = 'd1020;
    mem[11596] = 'd0;
    mem[11597] = 'd0;
    mem[11598] = 'd0;
    mem[11599] = 'd824;
    mem[11600] = 'd0;
    mem[11601] = 'd1020;
    mem[11602] = 'd0;
    mem[11603] = 'd0;
    mem[11604] = 'd0;
    mem[11605] = 'd820;
    mem[11606] = 'd0;
    mem[11607] = 'd1020;
    mem[11608] = 'd0;
    mem[11609] = 'd0;
    mem[11610] = 'd0;
    mem[11611] = 'd812;
    mem[11612] = 'd0;
    mem[11613] = 'd1020;
    mem[11614] = 'd0;
    mem[11615] = 'd0;
    mem[11616] = 'd0;
    mem[11617] = 'd772;
    mem[11618] = 'd0;
    mem[11619] = 'd1000;
    mem[11620] = 'd0;
    mem[11621] = 'd0;
    mem[11622] = 'd0;
    mem[11623] = 'd436;
    mem[11624] = 'd0;
    mem[11625] = 'd680;
    mem[11626] = 'd0;
    mem[11627] = 'd0;
    mem[11628] = 'd0;
    mem[11629] = 'd544;
    mem[11630] = 'd0;
    mem[11631] = 'd760;
    mem[11632] = 'd0;
    mem[11633] = 'd0;
    mem[11634] = 'd0;
    mem[11635] = 'd772;
    mem[11636] = 'd0;
    mem[11637] = 'd1020;
    mem[11638] = 'd0;
    mem[11639] = 'd0;
    mem[11640] = 'd0;
    mem[11641] = 'd756;
    mem[11642] = 'd0;
    mem[11643] = 'd1020;
    mem[11644] = 'd0;
    mem[11645] = 'd0;
    mem[11646] = 'd0;
    mem[11647] = 'd736;
    mem[11648] = 'd0;
    mem[11649] = 'd1016;
    mem[11650] = 'd0;
    mem[11651] = 'd0;
    mem[11652] = 'd0;
    mem[11653] = 'd720;
    mem[11654] = 'd0;
    mem[11655] = 'd1012;
    mem[11656] = 'd0;
    mem[11657] = 'd0;
    mem[11658] = 'd0;
    mem[11659] = 'd684;
    mem[11660] = 'd0;
    mem[11661] = 'd1000;
    mem[11662] = 'd0;
    mem[11663] = 'd0;
    mem[11664] = 'd0;
    mem[11665] = 'd636;
    mem[11666] = 'd0;
    mem[11667] = 'd956;
    mem[11668] = 'd0;
    mem[11669] = 'd0;
    mem[11670] = 'd0;
    mem[11671] = 'd556;
    mem[11672] = 'd0;
    mem[11673] = 'd904;
    mem[11674] = 'd0;
    mem[11675] = 'd0;
    mem[11676] = 'd0;
    mem[11677] = 'd464;
    mem[11678] = 'd0;
    mem[11679] = 'd840;
    mem[11680] = 'd0;
    mem[11681] = 'd0;
    mem[11682] = 'd0;
    mem[11683] = 'd952;
    mem[11684] = 'd0;
    mem[11685] = 'd984;
    mem[11686] = 'd0;
    mem[11687] = 'd0;
    mem[11688] = 'd0;
    mem[11689] = 'd1020;
    mem[11690] = 'd0;
    mem[11691] = 'd1020;
    mem[11692] = 'd0;
    mem[11693] = 'd0;
    mem[11694] = 'd0;
    mem[11695] = 'd1020;
    mem[11696] = 'd0;
    mem[11697] = 'd1020;
    mem[11698] = 'd0;
    mem[11699] = 'd0;
    mem[11700] = 'd0;
    mem[11701] = 'd0;
    mem[11702] = 'd1020;
    mem[11703] = 'd0;
    mem[11704] = 'd1020;
    mem[11705] = 'd0;
    mem[11706] = 'd0;
    mem[11707] = 'd0;
    mem[11708] = 'd1020;
    mem[11709] = 'd0;
    mem[11710] = 'd1020;
    mem[11711] = 'd0;
    mem[11712] = 'd0;
    mem[11713] = 'd0;
    mem[11714] = 'd356;
    mem[11715] = 'd0;
    mem[11716] = 'd624;
    mem[11717] = 'd0;
    mem[11718] = 'd0;
    mem[11719] = 'd0;
    mem[11720] = 'd24;
    mem[11721] = 'd0;
    mem[11722] = 'd504;
    mem[11723] = 'd0;
    mem[11724] = 'd0;
    mem[11725] = 'd0;
    mem[11726] = 'd52;
    mem[11727] = 'd0;
    mem[11728] = 'd600;
    mem[11729] = 'd0;
    mem[11730] = 'd0;
    mem[11731] = 'd0;
    mem[11732] = 'd68;
    mem[11733] = 'd0;
    mem[11734] = 'd656;
    mem[11735] = 'd0;
    mem[11736] = 'd0;
    mem[11737] = 'd0;
    mem[11738] = 'd84;
    mem[11739] = 'd0;
    mem[11740] = 'd692;
    mem[11741] = 'd0;
    mem[11742] = 'd0;
    mem[11743] = 'd0;
    mem[11744] = 'd112;
    mem[11745] = 'd0;
    mem[11746] = 'd720;
    mem[11747] = 'd0;
    mem[11748] = 'd0;
    mem[11749] = 'd0;
    mem[11750] = 'd160;
    mem[11751] = 'd0;
    mem[11752] = 'd740;
    mem[11753] = 'd0;
    mem[11754] = 'd0;
    mem[11755] = 'd0;
    mem[11756] = 'd192;
    mem[11757] = 'd0;
    mem[11758] = 'd756;
    mem[11759] = 'd0;
    mem[11760] = 'd0;
    mem[11761] = 'd0;
    mem[11762] = 'd224;
    mem[11763] = 'd0;
    mem[11764] = 'd736;
    mem[11765] = 'd0;
    mem[11766] = 'd0;
    mem[11767] = 'd0;
    mem[11768] = 'd44;
    mem[11769] = 'd0;
    mem[11770] = 'd288;
    mem[11771] = 'd0;
    mem[11772] = 'd0;
    mem[11773] = 'd0;
    mem[11774] = 'd44;
    mem[11775] = 'd0;
    mem[11776] = 'd332;
    mem[11777] = 'd0;
    mem[11778] = 'd0;
    mem[11779] = 'd0;
    mem[11780] = 'd128;
    mem[11781] = 'd0;
    mem[11782] = 'd572;
    mem[11783] = 'd0;
    mem[11784] = 'd0;
    mem[11785] = 'd0;
    mem[11786] = 'd204;
    mem[11787] = 'd0;
    mem[11788] = 'd764;
    mem[11789] = 'd0;
    mem[11790] = 'd0;
    mem[11791] = 'd0;
    mem[11792] = 'd224;
    mem[11793] = 'd0;
    mem[11794] = 'd804;
    mem[11795] = 'd0;
    mem[11796] = 'd0;
    mem[11797] = 'd0;
    mem[11798] = 'd228;
    mem[11799] = 'd0;
    mem[11800] = 'd812;
    mem[11801] = 'd0;
    mem[11802] = 'd0;
    mem[11803] = 'd0;
    mem[11804] = 'd228;
    mem[11805] = 'd0;
    mem[11806] = 'd812;
    mem[11807] = 'd0;
    mem[11808] = 'd0;
    mem[11809] = 'd0;
    mem[11810] = 'd228;
    mem[11811] = 'd0;
    mem[11812] = 'd816;
    mem[11813] = 'd0;
    mem[11814] = 'd0;
    mem[11815] = 'd0;
    mem[11816] = 'd228;
    mem[11817] = 'd0;
    mem[11818] = 'd816;
    mem[11819] = 'd0;
    mem[11820] = 'd0;
    mem[11821] = 'd0;
    mem[11822] = 'd228;
    mem[11823] = 'd0;
    mem[11824] = 'd812;
    mem[11825] = 'd0;
    mem[11826] = 'd0;
    mem[11827] = 'd0;
    mem[11828] = 'd224;
    mem[11829] = 'd0;
    mem[11830] = 'd808;
    mem[11831] = 'd0;
    mem[11832] = 'd0;
    mem[11833] = 'd0;
    mem[11834] = 'd220;
    mem[11835] = 'd0;
    mem[11836] = 'd796;
    mem[11837] = 'd0;
    mem[11838] = 'd0;
    mem[11839] = 'd0;
    mem[11840] = 'd192;
    mem[11841] = 'd0;
    mem[11842] = 'd736;
    mem[11843] = 'd0;
    mem[11844] = 'd0;
    mem[11845] = 'd0;
    mem[11846] = 'd116;
    mem[11847] = 'd0;
    mem[11848] = 'd532;
    mem[11849] = 'd0;
    mem[11850] = 'd0;
    mem[11851] = 'd0;
    mem[11852] = 'd36;
    mem[11853] = 'd0;
    mem[11854] = 'd300;
    mem[11855] = 'd0;
    mem[11856] = 'd0;
    mem[11857] = 'd0;
    mem[11858] = 'd64;
    mem[11859] = 'd0;
    mem[11860] = 'd328;
    mem[11861] = 'd0;
    mem[11862] = 'd0;
    mem[11863] = 'd0;
    mem[11864] = 'd236;
    mem[11865] = 'd0;
    mem[11866] = 'd772;
    mem[11867] = 'd0;
    mem[11868] = 'd0;
    mem[11869] = 'd0;
    mem[11870] = 'd196;
    mem[11871] = 'd0;
    mem[11872] = 'd752;
    mem[11873] = 'd0;
    mem[11874] = 'd0;
    mem[11875] = 'd0;
    mem[11876] = 'd160;
    mem[11877] = 'd0;
    mem[11878] = 'd740;
    mem[11879] = 'd0;
    mem[11880] = 'd0;
    mem[11881] = 'd0;
    mem[11882] = 'd116;
    mem[11883] = 'd0;
    mem[11884] = 'd724;
    mem[11885] = 'd0;
    mem[11886] = 'd0;
    mem[11887] = 'd0;
    mem[11888] = 'd84;
    mem[11889] = 'd0;
    mem[11890] = 'd696;
    mem[11891] = 'd0;
    mem[11892] = 'd0;
    mem[11893] = 'd0;
    mem[11894] = 'd72;
    mem[11895] = 'd0;
    mem[11896] = 'd660;
    mem[11897] = 'd0;
    mem[11898] = 'd0;
    mem[11899] = 'd0;
    mem[11900] = 'd56;
    mem[11901] = 'd0;
    mem[11902] = 'd604;
    mem[11903] = 'd0;
    mem[11904] = 'd0;
    mem[11905] = 'd0;
    mem[11906] = 'd28;
    mem[11907] = 'd0;
    mem[11908] = 'd508;
    mem[11909] = 'd0;
    mem[11910] = 'd0;
    mem[11911] = 'd0;
    mem[11912] = 'd292;
    mem[11913] = 'd0;
    mem[11914] = 'd584;
    mem[11915] = 'd0;
    mem[11916] = 'd0;
    mem[11917] = 'd0;
    mem[11918] = 'd1020;
    mem[11919] = 'd0;
    mem[11920] = 'd1020;
    mem[11921] = 'd0;
    mem[11922] = 'd0;
    mem[11923] = 'd0;
    mem[11924] = 'd1020;
    mem[11925] = 'd0;
    mem[11926] = 'd1020;
    mem[11927] = 'd0;
    mem[11928] = 'd0;
    mem[11929] = 'd0;
    mem[11930] = 'd1020;
    mem[11931] = 'd0;
    mem[11932] = 'd1020;
    mem[11933] = 'd0;
    mem[11934] = 'd0;
    mem[11935] = 'd1020;
    mem[11936] = 'd0;
    mem[11937] = 'd1020;
    mem[11938] = 'd0;
    mem[11939] = 'd0;
    mem[11940] = 'd0;
    mem[11941] = 'd1020;
    mem[11942] = 'd0;
    mem[11943] = 'd1020;
    mem[11944] = 'd0;
    mem[11945] = 'd0;
    mem[11946] = 'd0;
    mem[11947] = 'd624;
    mem[11948] = 'd0;
    mem[11949] = 'd876;
    mem[11950] = 'd0;
    mem[11951] = 'd0;
    mem[11952] = 'd0;
    mem[11953] = 'd504;
    mem[11954] = 'd0;
    mem[11955] = 'd860;
    mem[11956] = 'd0;
    mem[11957] = 'd0;
    mem[11958] = 'd0;
    mem[11959] = 'd600;
    mem[11960] = 'd0;
    mem[11961] = 'd924;
    mem[11962] = 'd0;
    mem[11963] = 'd0;
    mem[11964] = 'd0;
    mem[11965] = 'd656;
    mem[11966] = 'd0;
    mem[11967] = 'd972;
    mem[11968] = 'd0;
    mem[11969] = 'd0;
    mem[11970] = 'd0;
    mem[11971] = 'd692;
    mem[11972] = 'd0;
    mem[11973] = 'd1004;
    mem[11974] = 'd0;
    mem[11975] = 'd0;
    mem[11976] = 'd0;
    mem[11977] = 'd720;
    mem[11978] = 'd0;
    mem[11979] = 'd1016;
    mem[11980] = 'd0;
    mem[11981] = 'd0;
    mem[11982] = 'd0;
    mem[11983] = 'd740;
    mem[11984] = 'd0;
    mem[11985] = 'd1016;
    mem[11986] = 'd0;
    mem[11987] = 'd0;
    mem[11988] = 'd0;
    mem[11989] = 'd756;
    mem[11990] = 'd0;
    mem[11991] = 'd1020;
    mem[11992] = 'd0;
    mem[11993] = 'd0;
    mem[11994] = 'd0;
    mem[11995] = 'd736;
    mem[11996] = 'd0;
    mem[11997] = 'd948;
    mem[11998] = 'd0;
    mem[11999] = 'd0;
    mem[12000] = 'd0;
    mem[12001] = 'd288;
    mem[12002] = 'd0;
    mem[12003] = 'd500;
    mem[12004] = 'd0;
    mem[12005] = 'd0;
    mem[12006] = 'd0;
    mem[12007] = 'd332;
    mem[12008] = 'd0;
    mem[12009] = 'd564;
    mem[12010] = 'd0;
    mem[12011] = 'd0;
    mem[12012] = 'd0;
    mem[12013] = 'd572;
    mem[12014] = 'd0;
    mem[12015] = 'd820;
    mem[12016] = 'd0;
    mem[12017] = 'd0;
    mem[12018] = 'd0;
    mem[12019] = 'd764;
    mem[12020] = 'd0;
    mem[12021] = 'd1000;
    mem[12022] = 'd0;
    mem[12023] = 'd0;
    mem[12024] = 'd0;
    mem[12025] = 'd804;
    mem[12026] = 'd0;
    mem[12027] = 'd1016;
    mem[12028] = 'd0;
    mem[12029] = 'd0;
    mem[12030] = 'd0;
    mem[12031] = 'd812;
    mem[12032] = 'd0;
    mem[12033] = 'd1020;
    mem[12034] = 'd0;
    mem[12035] = 'd0;
    mem[12036] = 'd0;
    mem[12037] = 'd812;
    mem[12038] = 'd0;
    mem[12039] = 'd1020;
    mem[12040] = 'd0;
    mem[12041] = 'd0;
    mem[12042] = 'd0;
    mem[12043] = 'd816;
    mem[12044] = 'd0;
    mem[12045] = 'd1020;
    mem[12046] = 'd0;
    mem[12047] = 'd0;
    mem[12048] = 'd0;
    mem[12049] = 'd816;
    mem[12050] = 'd0;
    mem[12051] = 'd1020;
    mem[12052] = 'd0;
    mem[12053] = 'd0;
    mem[12054] = 'd0;
    mem[12055] = 'd812;
    mem[12056] = 'd0;
    mem[12057] = 'd1020;
    mem[12058] = 'd0;
    mem[12059] = 'd0;
    mem[12060] = 'd0;
    mem[12061] = 'd808;
    mem[12062] = 'd0;
    mem[12063] = 'd1020;
    mem[12064] = 'd0;
    mem[12065] = 'd0;
    mem[12066] = 'd0;
    mem[12067] = 'd796;
    mem[12068] = 'd0;
    mem[12069] = 'd1016;
    mem[12070] = 'd0;
    mem[12071] = 'd0;
    mem[12072] = 'd0;
    mem[12073] = 'd736;
    mem[12074] = 'd0;
    mem[12075] = 'd972;
    mem[12076] = 'd0;
    mem[12077] = 'd0;
    mem[12078] = 'd0;
    mem[12079] = 'd532;
    mem[12080] = 'd0;
    mem[12081] = 'd780;
    mem[12082] = 'd0;
    mem[12083] = 'd0;
    mem[12084] = 'd0;
    mem[12085] = 'd300;
    mem[12086] = 'd0;
    mem[12087] = 'd528;
    mem[12088] = 'd0;
    mem[12089] = 'd0;
    mem[12090] = 'd0;
    mem[12091] = 'd328;
    mem[12092] = 'd0;
    mem[12093] = 'd528;
    mem[12094] = 'd0;
    mem[12095] = 'd0;
    mem[12096] = 'd0;
    mem[12097] = 'd772;
    mem[12098] = 'd0;
    mem[12099] = 'd988;
    mem[12100] = 'd0;
    mem[12101] = 'd0;
    mem[12102] = 'd0;
    mem[12103] = 'd752;
    mem[12104] = 'd0;
    mem[12105] = 'd1020;
    mem[12106] = 'd0;
    mem[12107] = 'd0;
    mem[12108] = 'd0;
    mem[12109] = 'd740;
    mem[12110] = 'd0;
    mem[12111] = 'd1016;
    mem[12112] = 'd0;
    mem[12113] = 'd0;
    mem[12114] = 'd0;
    mem[12115] = 'd724;
    mem[12116] = 'd0;
    mem[12117] = 'd1016;
    mem[12118] = 'd0;
    mem[12119] = 'd0;
    mem[12120] = 'd0;
    mem[12121] = 'd696;
    mem[12122] = 'd0;
    mem[12123] = 'd1004;
    mem[12124] = 'd0;
    mem[12125] = 'd0;
    mem[12126] = 'd0;
    mem[12127] = 'd660;
    mem[12128] = 'd0;
    mem[12129] = 'd972;
    mem[12130] = 'd0;
    mem[12131] = 'd0;
    mem[12132] = 'd0;
    mem[12133] = 'd604;
    mem[12134] = 'd0;
    mem[12135] = 'd928;
    mem[12136] = 'd0;
    mem[12137] = 'd0;
    mem[12138] = 'd0;
    mem[12139] = 'd508;
    mem[12140] = 'd0;
    mem[12141] = 'd868;
    mem[12142] = 'd0;
    mem[12143] = 'd0;
    mem[12144] = 'd0;
    mem[12145] = 'd584;
    mem[12146] = 'd0;
    mem[12147] = 'd864;
    mem[12148] = 'd0;
    mem[12149] = 'd0;
    mem[12150] = 'd0;
    mem[12151] = 'd1020;
    mem[12152] = 'd0;
    mem[12153] = 'd1020;
    mem[12154] = 'd0;
    mem[12155] = 'd0;
    mem[12156] = 'd0;
    mem[12157] = 'd1020;
    mem[12158] = 'd0;
    mem[12159] = 'd1020;
    mem[12160] = 'd0;
    mem[12161] = 'd0;
    mem[12162] = 'd0;
    mem[12163] = 'd1020;
    mem[12164] = 'd0;
    mem[12165] = 'd1020;
    mem[12166] = 'd0;
    mem[12167] = 'd0;
    mem[12168] = 'd0;
    mem[12169] = 'd0;
    mem[12170] = 'd1020;
    mem[12171] = 'd0;
    mem[12172] = 'd1020;
    mem[12173] = 'd0;
    mem[12174] = 'd0;
    mem[12175] = 'd0;
    mem[12176] = 'd1020;
    mem[12177] = 'd0;
    mem[12178] = 'd1020;
    mem[12179] = 'd0;
    mem[12180] = 'd0;
    mem[12181] = 'd0;
    mem[12182] = 'd792;
    mem[12183] = 'd0;
    mem[12184] = 'd876;
    mem[12185] = 'd0;
    mem[12186] = 'd0;
    mem[12187] = 'd0;
    mem[12188] = 'd12;
    mem[12189] = 'd0;
    mem[12190] = 'd456;
    mem[12191] = 'd0;
    mem[12192] = 'd0;
    mem[12193] = 'd0;
    mem[12194] = 'd40;
    mem[12195] = 'd0;
    mem[12196] = 'd556;
    mem[12197] = 'd0;
    mem[12198] = 'd0;
    mem[12199] = 'd0;
    mem[12200] = 'd64;
    mem[12201] = 'd0;
    mem[12202] = 'd624;
    mem[12203] = 'd0;
    mem[12204] = 'd0;
    mem[12205] = 'd0;
    mem[12206] = 'd80;
    mem[12207] = 'd0;
    mem[12208] = 'd668;
    mem[12209] = 'd0;
    mem[12210] = 'd0;
    mem[12211] = 'd0;
    mem[12212] = 'd88;
    mem[12213] = 'd0;
    mem[12214] = 'd700;
    mem[12215] = 'd0;
    mem[12216] = 'd0;
    mem[12217] = 'd0;
    mem[12218] = 'd116;
    mem[12219] = 'd0;
    mem[12220] = 'd716;
    mem[12221] = 'd0;
    mem[12222] = 'd0;
    mem[12223] = 'd0;
    mem[12224] = 'd156;
    mem[12225] = 'd0;
    mem[12226] = 'd736;
    mem[12227] = 'd0;
    mem[12228] = 'd0;
    mem[12229] = 'd0;
    mem[12230] = 'd192;
    mem[12231] = 'd0;
    mem[12232] = 'd752;
    mem[12233] = 'd0;
    mem[12234] = 'd0;
    mem[12235] = 'd0;
    mem[12236] = 'd216;
    mem[12237] = 'd0;
    mem[12238] = 'd712;
    mem[12239] = 'd0;
    mem[12240] = 'd0;
    mem[12241] = 'd0;
    mem[12242] = 'd48;
    mem[12243] = 'd0;
    mem[12244] = 'd332;
    mem[12245] = 'd0;
    mem[12246] = 'd0;
    mem[12247] = 'd0;
    mem[12248] = 'd20;
    mem[12249] = 'd0;
    mem[12250] = 'd252;
    mem[12251] = 'd0;
    mem[12252] = 'd0;
    mem[12253] = 'd0;
    mem[12254] = 'd32;
    mem[12255] = 'd0;
    mem[12256] = 'd288;
    mem[12257] = 'd0;
    mem[12258] = 'd0;
    mem[12259] = 'd0;
    mem[12260] = 'd76;
    mem[12261] = 'd0;
    mem[12262] = 'd420;
    mem[12263] = 'd0;
    mem[12264] = 'd0;
    mem[12265] = 'd0;
    mem[12266] = 'd120;
    mem[12267] = 'd0;
    mem[12268] = 'd548;
    mem[12269] = 'd0;
    mem[12270] = 'd0;
    mem[12271] = 'd0;
    mem[12272] = 'd152;
    mem[12273] = 'd0;
    mem[12274] = 'd640;
    mem[12275] = 'd0;
    mem[12276] = 'd0;
    mem[12277] = 'd0;
    mem[12278] = 'd168;
    mem[12279] = 'd0;
    mem[12280] = 'd676;
    mem[12281] = 'd0;
    mem[12282] = 'd0;
    mem[12283] = 'd0;
    mem[12284] = 'd164;
    mem[12285] = 'd0;
    mem[12286] = 'd672;
    mem[12287] = 'd0;
    mem[12288] = 'd0;
    mem[12289] = 'd0;
    mem[12290] = 'd152;
    mem[12291] = 'd0;
    mem[12292] = 'd628;
    mem[12293] = 'd0;
    mem[12294] = 'd0;
    mem[12295] = 'd0;
    mem[12296] = 'd116;
    mem[12297] = 'd0;
    mem[12298] = 'd536;
    mem[12299] = 'd0;
    mem[12300] = 'd0;
    mem[12301] = 'd0;
    mem[12302] = 'd72;
    mem[12303] = 'd0;
    mem[12304] = 'd404;
    mem[12305] = 'd0;
    mem[12306] = 'd0;
    mem[12307] = 'd0;
    mem[12308] = 'd32;
    mem[12309] = 'd0;
    mem[12310] = 'd288;
    mem[12311] = 'd0;
    mem[12312] = 'd0;
    mem[12313] = 'd0;
    mem[12314] = 'd16;
    mem[12315] = 'd0;
    mem[12316] = 'd256;
    mem[12317] = 'd0;
    mem[12318] = 'd0;
    mem[12319] = 'd0;
    mem[12320] = 'd68;
    mem[12321] = 'd0;
    mem[12322] = 'd372;
    mem[12323] = 'd0;
    mem[12324] = 'd0;
    mem[12325] = 'd0;
    mem[12326] = 'd232;
    mem[12327] = 'd0;
    mem[12328] = 'd752;
    mem[12329] = 'd0;
    mem[12330] = 'd0;
    mem[12331] = 'd0;
    mem[12332] = 'd188;
    mem[12333] = 'd0;
    mem[12334] = 'd752;
    mem[12335] = 'd0;
    mem[12336] = 'd0;
    mem[12337] = 'd0;
    mem[12338] = 'd156;
    mem[12339] = 'd0;
    mem[12340] = 'd736;
    mem[12341] = 'd0;
    mem[12342] = 'd0;
    mem[12343] = 'd0;
    mem[12344] = 'd116;
    mem[12345] = 'd0;
    mem[12346] = 'd720;
    mem[12347] = 'd0;
    mem[12348] = 'd0;
    mem[12349] = 'd0;
    mem[12350] = 'd92;
    mem[12351] = 'd0;
    mem[12352] = 'd696;
    mem[12353] = 'd0;
    mem[12354] = 'd0;
    mem[12355] = 'd0;
    mem[12356] = 'd80;
    mem[12357] = 'd0;
    mem[12358] = 'd668;
    mem[12359] = 'd0;
    mem[12360] = 'd0;
    mem[12361] = 'd0;
    mem[12362] = 'd68;
    mem[12363] = 'd0;
    mem[12364] = 'd628;
    mem[12365] = 'd0;
    mem[12366] = 'd0;
    mem[12367] = 'd0;
    mem[12368] = 'd44;
    mem[12369] = 'd0;
    mem[12370] = 'd556;
    mem[12371] = 'd0;
    mem[12372] = 'd0;
    mem[12373] = 'd0;
    mem[12374] = 'd20;
    mem[12375] = 'd0;
    mem[12376] = 'd464;
    mem[12377] = 'd0;
    mem[12378] = 'd0;
    mem[12379] = 'd0;
    mem[12380] = 'd744;
    mem[12381] = 'd0;
    mem[12382] = 'd848;
    mem[12383] = 'd0;
    mem[12384] = 'd0;
    mem[12385] = 'd0;
    mem[12386] = 'd1020;
    mem[12387] = 'd0;
    mem[12388] = 'd1020;
    mem[12389] = 'd0;
    mem[12390] = 'd0;
    mem[12391] = 'd0;
    mem[12392] = 'd1020;
    mem[12393] = 'd0;
    mem[12394] = 'd1020;
    mem[12395] = 'd0;
    mem[12396] = 'd0;
    mem[12397] = 'd0;
    mem[12398] = 'd1020;
    mem[12399] = 'd0;
    mem[12400] = 'd1020;
    mem[12401] = 'd0;
    mem[12402] = 'd0;
    mem[12403] = 'd1020;
    mem[12404] = 'd0;
    mem[12405] = 'd1020;
    mem[12406] = 'd0;
    mem[12407] = 'd0;
    mem[12408] = 'd0;
    mem[12409] = 'd1020;
    mem[12410] = 'd0;
    mem[12411] = 'd1020;
    mem[12412] = 'd0;
    mem[12413] = 'd0;
    mem[12414] = 'd0;
    mem[12415] = 'd876;
    mem[12416] = 'd0;
    mem[12417] = 'd956;
    mem[12418] = 'd0;
    mem[12419] = 'd0;
    mem[12420] = 'd0;
    mem[12421] = 'd456;
    mem[12422] = 'd0;
    mem[12423] = 'd836;
    mem[12424] = 'd0;
    mem[12425] = 'd0;
    mem[12426] = 'd0;
    mem[12427] = 'd556;
    mem[12428] = 'd0;
    mem[12429] = 'd892;
    mem[12430] = 'd0;
    mem[12431] = 'd0;
    mem[12432] = 'd0;
    mem[12433] = 'd624;
    mem[12434] = 'd0;
    mem[12435] = 'd940;
    mem[12436] = 'd0;
    mem[12437] = 'd0;
    mem[12438] = 'd0;
    mem[12439] = 'd668;
    mem[12440] = 'd0;
    mem[12441] = 'd980;
    mem[12442] = 'd0;
    mem[12443] = 'd0;
    mem[12444] = 'd0;
    mem[12445] = 'd700;
    mem[12446] = 'd0;
    mem[12447] = 'd1008;
    mem[12448] = 'd0;
    mem[12449] = 'd0;
    mem[12450] = 'd0;
    mem[12451] = 'd716;
    mem[12452] = 'd0;
    mem[12453] = 'd1016;
    mem[12454] = 'd0;
    mem[12455] = 'd0;
    mem[12456] = 'd0;
    mem[12457] = 'd736;
    mem[12458] = 'd0;
    mem[12459] = 'd1020;
    mem[12460] = 'd0;
    mem[12461] = 'd0;
    mem[12462] = 'd0;
    mem[12463] = 'd752;
    mem[12464] = 'd0;
    mem[12465] = 'd1020;
    mem[12466] = 'd0;
    mem[12467] = 'd0;
    mem[12468] = 'd0;
    mem[12469] = 'd712;
    mem[12470] = 'd0;
    mem[12471] = 'd912;
    mem[12472] = 'd0;
    mem[12473] = 'd0;
    mem[12474] = 'd0;
    mem[12475] = 'd332;
    mem[12476] = 'd0;
    mem[12477] = 'd552;
    mem[12478] = 'd0;
    mem[12479] = 'd0;
    mem[12480] = 'd0;
    mem[12481] = 'd252;
    mem[12482] = 'd0;
    mem[12483] = 'd476;
    mem[12484] = 'd0;
    mem[12485] = 'd0;
    mem[12486] = 'd0;
    mem[12487] = 'd288;
    mem[12488] = 'd0;
    mem[12489] = 'd520;
    mem[12490] = 'd0;
    mem[12491] = 'd0;
    mem[12492] = 'd0;
    mem[12493] = 'd420;
    mem[12494] = 'd0;
    mem[12495] = 'd668;
    mem[12496] = 'd0;
    mem[12497] = 'd0;
    mem[12498] = 'd0;
    mem[12499] = 'd548;
    mem[12500] = 'd0;
    mem[12501] = 'd804;
    mem[12502] = 'd0;
    mem[12503] = 'd0;
    mem[12504] = 'd0;
    mem[12505] = 'd640;
    mem[12506] = 'd0;
    mem[12507] = 'd892;
    mem[12508] = 'd0;
    mem[12509] = 'd0;
    mem[12510] = 'd0;
    mem[12511] = 'd676;
    mem[12512] = 'd0;
    mem[12513] = 'd928;
    mem[12514] = 'd0;
    mem[12515] = 'd0;
    mem[12516] = 'd0;
    mem[12517] = 'd672;
    mem[12518] = 'd0;
    mem[12519] = 'd924;
    mem[12520] = 'd0;
    mem[12521] = 'd0;
    mem[12522] = 'd0;
    mem[12523] = 'd628;
    mem[12524] = 'd0;
    mem[12525] = 'd880;
    mem[12526] = 'd0;
    mem[12527] = 'd0;
    mem[12528] = 'd0;
    mem[12529] = 'd536;
    mem[12530] = 'd0;
    mem[12531] = 'd788;
    mem[12532] = 'd0;
    mem[12533] = 'd0;
    mem[12534] = 'd0;
    mem[12535] = 'd404;
    mem[12536] = 'd0;
    mem[12537] = 'd652;
    mem[12538] = 'd0;
    mem[12539] = 'd0;
    mem[12540] = 'd0;
    mem[12541] = 'd288;
    mem[12542] = 'd0;
    mem[12543] = 'd516;
    mem[12544] = 'd0;
    mem[12545] = 'd0;
    mem[12546] = 'd0;
    mem[12547] = 'd256;
    mem[12548] = 'd0;
    mem[12549] = 'd480;
    mem[12550] = 'd0;
    mem[12551] = 'd0;
    mem[12552] = 'd0;
    mem[12553] = 'd372;
    mem[12554] = 'd0;
    mem[12555] = 'd584;
    mem[12556] = 'd0;
    mem[12557] = 'd0;
    mem[12558] = 'd0;
    mem[12559] = 'd752;
    mem[12560] = 'd0;
    mem[12561] = 'd956;
    mem[12562] = 'd0;
    mem[12563] = 'd0;
    mem[12564] = 'd0;
    mem[12565] = 'd752;
    mem[12566] = 'd0;
    mem[12567] = 'd1020;
    mem[12568] = 'd0;
    mem[12569] = 'd0;
    mem[12570] = 'd0;
    mem[12571] = 'd736;
    mem[12572] = 'd0;
    mem[12573] = 'd1020;
    mem[12574] = 'd0;
    mem[12575] = 'd0;
    mem[12576] = 'd0;
    mem[12577] = 'd720;
    mem[12578] = 'd0;
    mem[12579] = 'd1016;
    mem[12580] = 'd0;
    mem[12581] = 'd0;
    mem[12582] = 'd0;
    mem[12583] = 'd696;
    mem[12584] = 'd0;
    mem[12585] = 'd1008;
    mem[12586] = 'd0;
    mem[12587] = 'd0;
    mem[12588] = 'd0;
    mem[12589] = 'd668;
    mem[12590] = 'd0;
    mem[12591] = 'd980;
    mem[12592] = 'd0;
    mem[12593] = 'd0;
    mem[12594] = 'd0;
    mem[12595] = 'd628;
    mem[12596] = 'd0;
    mem[12597] = 'd948;
    mem[12598] = 'd0;
    mem[12599] = 'd0;
    mem[12600] = 'd0;
    mem[12601] = 'd556;
    mem[12602] = 'd0;
    mem[12603] = 'd892;
    mem[12604] = 'd0;
    mem[12605] = 'd0;
    mem[12606] = 'd0;
    mem[12607] = 'd464;
    mem[12608] = 'd0;
    mem[12609] = 'd836;
    mem[12610] = 'd0;
    mem[12611] = 'd0;
    mem[12612] = 'd0;
    mem[12613] = 'd848;
    mem[12614] = 'd0;
    mem[12615] = 'd952;
    mem[12616] = 'd0;
    mem[12617] = 'd0;
    mem[12618] = 'd0;
    mem[12619] = 'd1020;
    mem[12620] = 'd0;
    mem[12621] = 'd1020;
    mem[12622] = 'd0;
    mem[12623] = 'd0;
    mem[12624] = 'd0;
    mem[12625] = 'd1020;
    mem[12626] = 'd0;
    mem[12627] = 'd1020;
    mem[12628] = 'd0;
    mem[12629] = 'd0;
    mem[12630] = 'd0;
    mem[12631] = 'd1020;
    mem[12632] = 'd0;
    mem[12633] = 'd1020;
    mem[12634] = 'd0;
    mem[12635] = 'd0;
    mem[12636] = 'd0;
    mem[12637] = 'd0;
    mem[12638] = 'd1020;
    mem[12639] = 'd0;
    mem[12640] = 'd1020;
    mem[12641] = 'd0;
    mem[12642] = 'd0;
    mem[12643] = 'd0;
    mem[12644] = 'd1020;
    mem[12645] = 'd0;
    mem[12646] = 'd1020;
    mem[12647] = 'd0;
    mem[12648] = 'd0;
    mem[12649] = 'd0;
    mem[12650] = 'd1020;
    mem[12651] = 'd0;
    mem[12652] = 'd1020;
    mem[12653] = 'd0;
    mem[12654] = 'd0;
    mem[12655] = 'd0;
    mem[12656] = 'd280;
    mem[12657] = 'd0;
    mem[12658] = 'd576;
    mem[12659] = 'd0;
    mem[12660] = 'd0;
    mem[12661] = 'd0;
    mem[12662] = 'd28;
    mem[12663] = 'd0;
    mem[12664] = 'd504;
    mem[12665] = 'd0;
    mem[12666] = 'd0;
    mem[12667] = 'd0;
    mem[12668] = 'd52;
    mem[12669] = 'd0;
    mem[12670] = 'd580;
    mem[12671] = 'd0;
    mem[12672] = 'd0;
    mem[12673] = 'd0;
    mem[12674] = 'd72;
    mem[12675] = 'd0;
    mem[12676] = 'd636;
    mem[12677] = 'd0;
    mem[12678] = 'd0;
    mem[12679] = 'd0;
    mem[12680] = 'd84;
    mem[12681] = 'd0;
    mem[12682] = 'd672;
    mem[12683] = 'd0;
    mem[12684] = 'd0;
    mem[12685] = 'd0;
    mem[12686] = 'd92;
    mem[12687] = 'd0;
    mem[12688] = 'd696;
    mem[12689] = 'd0;
    mem[12690] = 'd0;
    mem[12691] = 'd0;
    mem[12692] = 'd108;
    mem[12693] = 'd0;
    mem[12694] = 'd716;
    mem[12695] = 'd0;
    mem[12696] = 'd0;
    mem[12697] = 'd0;
    mem[12698] = 'd144;
    mem[12699] = 'd0;
    mem[12700] = 'd732;
    mem[12701] = 'd0;
    mem[12702] = 'd0;
    mem[12703] = 'd0;
    mem[12704] = 'd180;
    mem[12705] = 'd0;
    mem[12706] = 'd748;
    mem[12707] = 'd0;
    mem[12708] = 'd0;
    mem[12709] = 'd0;
    mem[12710] = 'd224;
    mem[12711] = 'd0;
    mem[12712] = 'd752;
    mem[12713] = 'd0;
    mem[12714] = 'd0;
    mem[12715] = 'd0;
    mem[12716] = 'd112;
    mem[12717] = 'd0;
    mem[12718] = 'd480;
    mem[12719] = 'd0;
    mem[12720] = 'd0;
    mem[12721] = 'd0;
    mem[12722] = 'd20;
    mem[12723] = 'd0;
    mem[12724] = 'd308;
    mem[12725] = 'd0;
    mem[12726] = 'd0;
    mem[12727] = 'd0;
    mem[12728] = 'd20;
    mem[12729] = 'd0;
    mem[12730] = 'd296;
    mem[12731] = 'd0;
    mem[12732] = 'd0;
    mem[12733] = 'd0;
    mem[12734] = 'd16;
    mem[12735] = 'd0;
    mem[12736] = 'd264;
    mem[12737] = 'd0;
    mem[12738] = 'd0;
    mem[12739] = 'd0;
    mem[12740] = 'd20;
    mem[12741] = 'd0;
    mem[12742] = 'd248;
    mem[12743] = 'd0;
    mem[12744] = 'd0;
    mem[12745] = 'd0;
    mem[12746] = 'd20;
    mem[12747] = 'd0;
    mem[12748] = 'd244;
    mem[12749] = 'd0;
    mem[12750] = 'd0;
    mem[12751] = 'd0;
    mem[12752] = 'd20;
    mem[12753] = 'd0;
    mem[12754] = 'd248;
    mem[12755] = 'd0;
    mem[12756] = 'd0;
    mem[12757] = 'd0;
    mem[12758] = 'd20;
    mem[12759] = 'd0;
    mem[12760] = 'd252;
    mem[12761] = 'd0;
    mem[12762] = 'd0;
    mem[12763] = 'd0;
    mem[12764] = 'd16;
    mem[12765] = 'd0;
    mem[12766] = 'd268;
    mem[12767] = 'd0;
    mem[12768] = 'd0;
    mem[12769] = 'd0;
    mem[12770] = 'd20;
    mem[12771] = 'd0;
    mem[12772] = 'd300;
    mem[12773] = 'd0;
    mem[12774] = 'd0;
    mem[12775] = 'd0;
    mem[12776] = 'd28;
    mem[12777] = 'd0;
    mem[12778] = 'd328;
    mem[12779] = 'd0;
    mem[12780] = 'd0;
    mem[12781] = 'd0;
    mem[12782] = 'd136;
    mem[12783] = 'd0;
    mem[12784] = 'd532;
    mem[12785] = 'd0;
    mem[12786] = 'd0;
    mem[12787] = 'd0;
    mem[12788] = 'd224;
    mem[12789] = 'd0;
    mem[12790] = 'd768;
    mem[12791] = 'd0;
    mem[12792] = 'd0;
    mem[12793] = 'd0;
    mem[12794] = 'd176;
    mem[12795] = 'd0;
    mem[12796] = 'd748;
    mem[12797] = 'd0;
    mem[12798] = 'd0;
    mem[12799] = 'd0;
    mem[12800] = 'd144;
    mem[12801] = 'd0;
    mem[12802] = 'd732;
    mem[12803] = 'd0;
    mem[12804] = 'd0;
    mem[12805] = 'd0;
    mem[12806] = 'd112;
    mem[12807] = 'd0;
    mem[12808] = 'd716;
    mem[12809] = 'd0;
    mem[12810] = 'd0;
    mem[12811] = 'd0;
    mem[12812] = 'd92;
    mem[12813] = 'd0;
    mem[12814] = 'd696;
    mem[12815] = 'd0;
    mem[12816] = 'd0;
    mem[12817] = 'd0;
    mem[12818] = 'd84;
    mem[12819] = 'd0;
    mem[12820] = 'd676;
    mem[12821] = 'd0;
    mem[12822] = 'd0;
    mem[12823] = 'd0;
    mem[12824] = 'd76;
    mem[12825] = 'd0;
    mem[12826] = 'd640;
    mem[12827] = 'd0;
    mem[12828] = 'd0;
    mem[12829] = 'd0;
    mem[12830] = 'd56;
    mem[12831] = 'd0;
    mem[12832] = 'd588;
    mem[12833] = 'd0;
    mem[12834] = 'd0;
    mem[12835] = 'd0;
    mem[12836] = 'd32;
    mem[12837] = 'd0;
    mem[12838] = 'd508;
    mem[12839] = 'd0;
    mem[12840] = 'd0;
    mem[12841] = 'd0;
    mem[12842] = 'd256;
    mem[12843] = 'd0;
    mem[12844] = 'd564;
    mem[12845] = 'd0;
    mem[12846] = 'd0;
    mem[12847] = 'd0;
    mem[12848] = 'd1008;
    mem[12849] = 'd0;
    mem[12850] = 'd1012;
    mem[12851] = 'd0;
    mem[12852] = 'd0;
    mem[12853] = 'd0;
    mem[12854] = 'd1020;
    mem[12855] = 'd0;
    mem[12856] = 'd1020;
    mem[12857] = 'd0;
    mem[12858] = 'd0;
    mem[12859] = 'd0;
    mem[12860] = 'd1020;
    mem[12861] = 'd0;
    mem[12862] = 'd1020;
    mem[12863] = 'd0;
    mem[12864] = 'd0;
    mem[12865] = 'd0;
    mem[12866] = 'd1020;
    mem[12867] = 'd0;
    mem[12868] = 'd1020;
    mem[12869] = 'd0;
    mem[12870] = 'd0;
    mem[12871] = 'd1020;
    mem[12872] = 'd0;
    mem[12873] = 'd1020;
    mem[12874] = 'd0;
    mem[12875] = 'd0;
    mem[12876] = 'd0;
    mem[12877] = 'd1020;
    mem[12878] = 'd0;
    mem[12879] = 'd1020;
    mem[12880] = 'd0;
    mem[12881] = 'd0;
    mem[12882] = 'd0;
    mem[12883] = 'd1020;
    mem[12884] = 'd0;
    mem[12885] = 'd1020;
    mem[12886] = 'd0;
    mem[12887] = 'd0;
    mem[12888] = 'd0;
    mem[12889] = 'd576;
    mem[12890] = 'd0;
    mem[12891] = 'd856;
    mem[12892] = 'd0;
    mem[12893] = 'd0;
    mem[12894] = 'd0;
    mem[12895] = 'd504;
    mem[12896] = 'd0;
    mem[12897] = 'd856;
    mem[12898] = 'd0;
    mem[12899] = 'd0;
    mem[12900] = 'd0;
    mem[12901] = 'd580;
    mem[12902] = 'd0;
    mem[12903] = 'd904;
    mem[12904] = 'd0;
    mem[12905] = 'd0;
    mem[12906] = 'd0;
    mem[12907] = 'd636;
    mem[12908] = 'd0;
    mem[12909] = 'd952;
    mem[12910] = 'd0;
    mem[12911] = 'd0;
    mem[12912] = 'd0;
    mem[12913] = 'd672;
    mem[12914] = 'd0;
    mem[12915] = 'd984;
    mem[12916] = 'd0;
    mem[12917] = 'd0;
    mem[12918] = 'd0;
    mem[12919] = 'd696;
    mem[12920] = 'd0;
    mem[12921] = 'd1004;
    mem[12922] = 'd0;
    mem[12923] = 'd0;
    mem[12924] = 'd0;
    mem[12925] = 'd716;
    mem[12926] = 'd0;
    mem[12927] = 'd1020;
    mem[12928] = 'd0;
    mem[12929] = 'd0;
    mem[12930] = 'd0;
    mem[12931] = 'd732;
    mem[12932] = 'd0;
    mem[12933] = 'd1020;
    mem[12934] = 'd0;
    mem[12935] = 'd0;
    mem[12936] = 'd0;
    mem[12937] = 'd748;
    mem[12938] = 'd0;
    mem[12939] = 'd1020;
    mem[12940] = 'd0;
    mem[12941] = 'd0;
    mem[12942] = 'd0;
    mem[12943] = 'd752;
    mem[12944] = 'd0;
    mem[12945] = 'd956;
    mem[12946] = 'd0;
    mem[12947] = 'd0;
    mem[12948] = 'd0;
    mem[12949] = 'd480;
    mem[12950] = 'd0;
    mem[12951] = 'd680;
    mem[12952] = 'd0;
    mem[12953] = 'd0;
    mem[12954] = 'd0;
    mem[12955] = 'd308;
    mem[12956] = 'd0;
    mem[12957] = 'd544;
    mem[12958] = 'd0;
    mem[12959] = 'd0;
    mem[12960] = 'd0;
    mem[12961] = 'd296;
    mem[12962] = 'd0;
    mem[12963] = 'd528;
    mem[12964] = 'd0;
    mem[12965] = 'd0;
    mem[12966] = 'd0;
    mem[12967] = 'd264;
    mem[12968] = 'd0;
    mem[12969] = 'd488;
    mem[12970] = 'd0;
    mem[12971] = 'd0;
    mem[12972] = 'd0;
    mem[12973] = 'd248;
    mem[12974] = 'd0;
    mem[12975] = 'd468;
    mem[12976] = 'd0;
    mem[12977] = 'd0;
    mem[12978] = 'd0;
    mem[12979] = 'd244;
    mem[12980] = 'd0;
    mem[12981] = 'd468;
    mem[12982] = 'd0;
    mem[12983] = 'd0;
    mem[12984] = 'd0;
    mem[12985] = 'd248;
    mem[12986] = 'd0;
    mem[12987] = 'd468;
    mem[12988] = 'd0;
    mem[12989] = 'd0;
    mem[12990] = 'd0;
    mem[12991] = 'd252;
    mem[12992] = 'd0;
    mem[12993] = 'd472;
    mem[12994] = 'd0;
    mem[12995] = 'd0;
    mem[12996] = 'd0;
    mem[12997] = 'd268;
    mem[12998] = 'd0;
    mem[12999] = 'd496;
    mem[13000] = 'd0;
    mem[13001] = 'd0;
    mem[13002] = 'd0;
    mem[13003] = 'd300;
    mem[13004] = 'd0;
    mem[13005] = 'd528;
    mem[13006] = 'd0;
    mem[13007] = 'd0;
    mem[13008] = 'd0;
    mem[13009] = 'd328;
    mem[13010] = 'd0;
    mem[13011] = 'd560;
    mem[13012] = 'd0;
    mem[13013] = 'd0;
    mem[13014] = 'd0;
    mem[13015] = 'd532;
    mem[13016] = 'd0;
    mem[13017] = 'd728;
    mem[13018] = 'd0;
    mem[13019] = 'd0;
    mem[13020] = 'd0;
    mem[13021] = 'd768;
    mem[13022] = 'd0;
    mem[13023] = 'd976;
    mem[13024] = 'd0;
    mem[13025] = 'd0;
    mem[13026] = 'd0;
    mem[13027] = 'd748;
    mem[13028] = 'd0;
    mem[13029] = 'd1020;
    mem[13030] = 'd0;
    mem[13031] = 'd0;
    mem[13032] = 'd0;
    mem[13033] = 'd732;
    mem[13034] = 'd0;
    mem[13035] = 'd1020;
    mem[13036] = 'd0;
    mem[13037] = 'd0;
    mem[13038] = 'd0;
    mem[13039] = 'd716;
    mem[13040] = 'd0;
    mem[13041] = 'd1020;
    mem[13042] = 'd0;
    mem[13043] = 'd0;
    mem[13044] = 'd0;
    mem[13045] = 'd696;
    mem[13046] = 'd0;
    mem[13047] = 'd1008;
    mem[13048] = 'd0;
    mem[13049] = 'd0;
    mem[13050] = 'd0;
    mem[13051] = 'd676;
    mem[13052] = 'd0;
    mem[13053] = 'd984;
    mem[13054] = 'd0;
    mem[13055] = 'd0;
    mem[13056] = 'd0;
    mem[13057] = 'd640;
    mem[13058] = 'd0;
    mem[13059] = 'd956;
    mem[13060] = 'd0;
    mem[13061] = 'd0;
    mem[13062] = 'd0;
    mem[13063] = 'd588;
    mem[13064] = 'd0;
    mem[13065] = 'd912;
    mem[13066] = 'd0;
    mem[13067] = 'd0;
    mem[13068] = 'd0;
    mem[13069] = 'd508;
    mem[13070] = 'd0;
    mem[13071] = 'd860;
    mem[13072] = 'd0;
    mem[13073] = 'd0;
    mem[13074] = 'd0;
    mem[13075] = 'd564;
    mem[13076] = 'd0;
    mem[13077] = 'd856;
    mem[13078] = 'd0;
    mem[13079] = 'd0;
    mem[13080] = 'd0;
    mem[13081] = 'd1012;
    mem[13082] = 'd0;
    mem[13083] = 'd1012;
    mem[13084] = 'd0;
    mem[13085] = 'd0;
    mem[13086] = 'd0;
    mem[13087] = 'd1020;
    mem[13088] = 'd0;
    mem[13089] = 'd1020;
    mem[13090] = 'd0;
    mem[13091] = 'd0;
    mem[13092] = 'd0;
    mem[13093] = 'd1020;
    mem[13094] = 'd0;
    mem[13095] = 'd1020;
    mem[13096] = 'd0;
    mem[13097] = 'd0;
    mem[13098] = 'd0;
    mem[13099] = 'd1020;
    mem[13100] = 'd0;
    mem[13101] = 'd1020;
    mem[13102] = 'd0;
    mem[13103] = 'd0;
    mem[13104] = 'd0;
    mem[13105] = 'd0;
    mem[13106] = 'd1020;
    mem[13107] = 'd0;
    mem[13108] = 'd1020;
    mem[13109] = 'd0;
    mem[13110] = 'd0;
    mem[13111] = 'd0;
    mem[13112] = 'd1020;
    mem[13113] = 'd0;
    mem[13114] = 'd1020;
    mem[13115] = 'd0;
    mem[13116] = 'd0;
    mem[13117] = 'd0;
    mem[13118] = 'd1020;
    mem[13119] = 'd0;
    mem[13120] = 'd1020;
    mem[13121] = 'd0;
    mem[13122] = 'd0;
    mem[13123] = 'd0;
    mem[13124] = 'd848;
    mem[13125] = 'd0;
    mem[13126] = 'd912;
    mem[13127] = 'd0;
    mem[13128] = 'd0;
    mem[13129] = 'd0;
    mem[13130] = 'd24;
    mem[13131] = 'd0;
    mem[13132] = 'd456;
    mem[13133] = 'd0;
    mem[13134] = 'd0;
    mem[13135] = 'd0;
    mem[13136] = 'd36;
    mem[13137] = 'd0;
    mem[13138] = 'd528;
    mem[13139] = 'd0;
    mem[13140] = 'd0;
    mem[13141] = 'd0;
    mem[13142] = 'd60;
    mem[13143] = 'd0;
    mem[13144] = 'd596;
    mem[13145] = 'd0;
    mem[13146] = 'd0;
    mem[13147] = 'd0;
    mem[13148] = 'd76;
    mem[13149] = 'd0;
    mem[13150] = 'd640;
    mem[13151] = 'd0;
    mem[13152] = 'd0;
    mem[13153] = 'd0;
    mem[13154] = 'd88;
    mem[13155] = 'd0;
    mem[13156] = 'd672;
    mem[13157] = 'd0;
    mem[13158] = 'd0;
    mem[13159] = 'd0;
    mem[13160] = 'd92;
    mem[13161] = 'd0;
    mem[13162] = 'd692;
    mem[13163] = 'd0;
    mem[13164] = 'd0;
    mem[13165] = 'd0;
    mem[13166] = 'd100;
    mem[13167] = 'd0;
    mem[13168] = 'd708;
    mem[13169] = 'd0;
    mem[13170] = 'd0;
    mem[13171] = 'd0;
    mem[13172] = 'd124;
    mem[13173] = 'd0;
    mem[13174] = 'd724;
    mem[13175] = 'd0;
    mem[13176] = 'd0;
    mem[13177] = 'd0;
    mem[13178] = 'd152;
    mem[13179] = 'd0;
    mem[13180] = 'd736;
    mem[13181] = 'd0;
    mem[13182] = 'd0;
    mem[13183] = 'd0;
    mem[13184] = 'd200;
    mem[13185] = 'd0;
    mem[13186] = 'd768;
    mem[13187] = 'd0;
    mem[13188] = 'd0;
    mem[13189] = 'd0;
    mem[13190] = 'd204;
    mem[13191] = 'd0;
    mem[13192] = 'd708;
    mem[13193] = 'd0;
    mem[13194] = 'd0;
    mem[13195] = 'd0;
    mem[13196] = 'd132;
    mem[13197] = 'd0;
    mem[13198] = 'd532;
    mem[13199] = 'd0;
    mem[13200] = 'd0;
    mem[13201] = 'd0;
    mem[13202] = 'd60;
    mem[13203] = 'd0;
    mem[13204] = 'd400;
    mem[13205] = 'd0;
    mem[13206] = 'd0;
    mem[13207] = 'd0;
    mem[13208] = 'd32;
    mem[13209] = 'd0;
    mem[13210] = 'd352;
    mem[13211] = 'd0;
    mem[13212] = 'd0;
    mem[13213] = 'd0;
    mem[13214] = 'd24;
    mem[13215] = 'd0;
    mem[13216] = 'd344;
    mem[13217] = 'd0;
    mem[13218] = 'd0;
    mem[13219] = 'd0;
    mem[13220] = 'd28;
    mem[13221] = 'd0;
    mem[13222] = 'd344;
    mem[13223] = 'd0;
    mem[13224] = 'd0;
    mem[13225] = 'd0;
    mem[13226] = 'd36;
    mem[13227] = 'd0;
    mem[13228] = 'd364;
    mem[13229] = 'd0;
    mem[13230] = 'd0;
    mem[13231] = 'd0;
    mem[13232] = 'd72;
    mem[13233] = 'd0;
    mem[13234] = 'd420;
    mem[13235] = 'd0;
    mem[13236] = 'd0;
    mem[13237] = 'd0;
    mem[13238] = 'd140;
    mem[13239] = 'd0;
    mem[13240] = 'd556;
    mem[13241] = 'd0;
    mem[13242] = 'd0;
    mem[13243] = 'd0;
    mem[13244] = 'd204;
    mem[13245] = 'd0;
    mem[13246] = 'd716;
    mem[13247] = 'd0;
    mem[13248] = 'd0;
    mem[13249] = 'd0;
    mem[13250] = 'd192;
    mem[13251] = 'd0;
    mem[13252] = 'd764;
    mem[13253] = 'd0;
    mem[13254] = 'd0;
    mem[13255] = 'd0;
    mem[13256] = 'd156;
    mem[13257] = 'd0;
    mem[13258] = 'd736;
    mem[13259] = 'd0;
    mem[13260] = 'd0;
    mem[13261] = 'd0;
    mem[13262] = 'd128;
    mem[13263] = 'd0;
    mem[13264] = 'd724;
    mem[13265] = 'd0;
    mem[13266] = 'd0;
    mem[13267] = 'd0;
    mem[13268] = 'd100;
    mem[13269] = 'd0;
    mem[13270] = 'd708;
    mem[13271] = 'd0;
    mem[13272] = 'd0;
    mem[13273] = 'd0;
    mem[13274] = 'd92;
    mem[13275] = 'd0;
    mem[13276] = 'd692;
    mem[13277] = 'd0;
    mem[13278] = 'd0;
    mem[13279] = 'd0;
    mem[13280] = 'd88;
    mem[13281] = 'd0;
    mem[13282] = 'd672;
    mem[13283] = 'd0;
    mem[13284] = 'd0;
    mem[13285] = 'd0;
    mem[13286] = 'd80;
    mem[13287] = 'd0;
    mem[13288] = 'd644;
    mem[13289] = 'd0;
    mem[13290] = 'd0;
    mem[13291] = 'd0;
    mem[13292] = 'd64;
    mem[13293] = 'd0;
    mem[13294] = 'd600;
    mem[13295] = 'd0;
    mem[13296] = 'd0;
    mem[13297] = 'd0;
    mem[13298] = 'd40;
    mem[13299] = 'd0;
    mem[13300] = 'd532;
    mem[13301] = 'd0;
    mem[13302] = 'd0;
    mem[13303] = 'd0;
    mem[13304] = 'd52;
    mem[13305] = 'd0;
    mem[13306] = 'd472;
    mem[13307] = 'd0;
    mem[13308] = 'd0;
    mem[13309] = 'd0;
    mem[13310] = 'd796;
    mem[13311] = 'd0;
    mem[13312] = 'd880;
    mem[13313] = 'd0;
    mem[13314] = 'd0;
    mem[13315] = 'd0;
    mem[13316] = 'd1020;
    mem[13317] = 'd0;
    mem[13318] = 'd1020;
    mem[13319] = 'd0;
    mem[13320] = 'd0;
    mem[13321] = 'd0;
    mem[13322] = 'd1020;
    mem[13323] = 'd0;
    mem[13324] = 'd1020;
    mem[13325] = 'd0;
    mem[13326] = 'd0;
    mem[13327] = 'd0;
    mem[13328] = 'd1020;
    mem[13329] = 'd0;
    mem[13330] = 'd1020;
    mem[13331] = 'd0;
    mem[13332] = 'd0;
    mem[13333] = 'd0;
    mem[13334] = 'd1020;
    mem[13335] = 'd0;
    mem[13336] = 'd1020;
    mem[13337] = 'd0;
    mem[13338] = 'd0;
    mem[13339] = 'd1020;
    mem[13340] = 'd0;
    mem[13341] = 'd1020;
    mem[13342] = 'd0;
    mem[13343] = 'd0;
    mem[13344] = 'd0;
    mem[13345] = 'd1020;
    mem[13346] = 'd0;
    mem[13347] = 'd1020;
    mem[13348] = 'd0;
    mem[13349] = 'd0;
    mem[13350] = 'd0;
    mem[13351] = 'd1020;
    mem[13352] = 'd0;
    mem[13353] = 'd1020;
    mem[13354] = 'd0;
    mem[13355] = 'd0;
    mem[13356] = 'd0;
    mem[13357] = 'd912;
    mem[13358] = 'd0;
    mem[13359] = 'd972;
    mem[13360] = 'd0;
    mem[13361] = 'd0;
    mem[13362] = 'd0;
    mem[13363] = 'd456;
    mem[13364] = 'd0;
    mem[13365] = 'd828;
    mem[13366] = 'd0;
    mem[13367] = 'd0;
    mem[13368] = 'd0;
    mem[13369] = 'd528;
    mem[13370] = 'd0;
    mem[13371] = 'd868;
    mem[13372] = 'd0;
    mem[13373] = 'd0;
    mem[13374] = 'd0;
    mem[13375] = 'd596;
    mem[13376] = 'd0;
    mem[13377] = 'd916;
    mem[13378] = 'd0;
    mem[13379] = 'd0;
    mem[13380] = 'd0;
    mem[13381] = 'd640;
    mem[13382] = 'd0;
    mem[13383] = 'd956;
    mem[13384] = 'd0;
    mem[13385] = 'd0;
    mem[13386] = 'd0;
    mem[13387] = 'd672;
    mem[13388] = 'd0;
    mem[13389] = 'd984;
    mem[13390] = 'd0;
    mem[13391] = 'd0;
    mem[13392] = 'd0;
    mem[13393] = 'd692;
    mem[13394] = 'd0;
    mem[13395] = 'd1004;
    mem[13396] = 'd0;
    mem[13397] = 'd0;
    mem[13398] = 'd0;
    mem[13399] = 'd708;
    mem[13400] = 'd0;
    mem[13401] = 'd1016;
    mem[13402] = 'd0;
    mem[13403] = 'd0;
    mem[13404] = 'd0;
    mem[13405] = 'd724;
    mem[13406] = 'd0;
    mem[13407] = 'd1020;
    mem[13408] = 'd0;
    mem[13409] = 'd0;
    mem[13410] = 'd0;
    mem[13411] = 'd736;
    mem[13412] = 'd0;
    mem[13413] = 'd1020;
    mem[13414] = 'd0;
    mem[13415] = 'd0;
    mem[13416] = 'd0;
    mem[13417] = 'd768;
    mem[13418] = 'd0;
    mem[13419] = 'd1016;
    mem[13420] = 'd0;
    mem[13421] = 'd0;
    mem[13422] = 'd0;
    mem[13423] = 'd708;
    mem[13424] = 'd0;
    mem[13425] = 'd896;
    mem[13426] = 'd0;
    mem[13427] = 'd0;
    mem[13428] = 'd0;
    mem[13429] = 'd532;
    mem[13430] = 'd0;
    mem[13431] = 'd728;
    mem[13432] = 'd0;
    mem[13433] = 'd0;
    mem[13434] = 'd0;
    mem[13435] = 'd400;
    mem[13436] = 'd0;
    mem[13437] = 'd624;
    mem[13438] = 'd0;
    mem[13439] = 'd0;
    mem[13440] = 'd0;
    mem[13441] = 'd352;
    mem[13442] = 'd0;
    mem[13443] = 'd584;
    mem[13444] = 'd0;
    mem[13445] = 'd0;
    mem[13446] = 'd0;
    mem[13447] = 'd344;
    mem[13448] = 'd0;
    mem[13449] = 'd576;
    mem[13450] = 'd0;
    mem[13451] = 'd0;
    mem[13452] = 'd0;
    mem[13453] = 'd344;
    mem[13454] = 'd0;
    mem[13455] = 'd580;
    mem[13456] = 'd0;
    mem[13457] = 'd0;
    mem[13458] = 'd0;
    mem[13459] = 'd364;
    mem[13460] = 'd0;
    mem[13461] = 'd596;
    mem[13462] = 'd0;
    mem[13463] = 'd0;
    mem[13464] = 'd0;
    mem[13465] = 'd420;
    mem[13466] = 'd0;
    mem[13467] = 'd640;
    mem[13468] = 'd0;
    mem[13469] = 'd0;
    mem[13470] = 'd0;
    mem[13471] = 'd556;
    mem[13472] = 'd0;
    mem[13473] = 'd752;
    mem[13474] = 'd0;
    mem[13475] = 'd0;
    mem[13476] = 'd0;
    mem[13477] = 'd716;
    mem[13478] = 'd0;
    mem[13479] = 'd916;
    mem[13480] = 'd0;
    mem[13481] = 'd0;
    mem[13482] = 'd0;
    mem[13483] = 'd764;
    mem[13484] = 'd0;
    mem[13485] = 'd1020;
    mem[13486] = 'd0;
    mem[13487] = 'd0;
    mem[13488] = 'd0;
    mem[13489] = 'd736;
    mem[13490] = 'd0;
    mem[13491] = 'd1020;
    mem[13492] = 'd0;
    mem[13493] = 'd0;
    mem[13494] = 'd0;
    mem[13495] = 'd724;
    mem[13496] = 'd0;
    mem[13497] = 'd1020;
    mem[13498] = 'd0;
    mem[13499] = 'd0;
    mem[13500] = 'd0;
    mem[13501] = 'd708;
    mem[13502] = 'd0;
    mem[13503] = 'd1016;
    mem[13504] = 'd0;
    mem[13505] = 'd0;
    mem[13506] = 'd0;
    mem[13507] = 'd692;
    mem[13508] = 'd0;
    mem[13509] = 'd1008;
    mem[13510] = 'd0;
    mem[13511] = 'd0;
    mem[13512] = 'd0;
    mem[13513] = 'd672;
    mem[13514] = 'd0;
    mem[13515] = 'd988;
    mem[13516] = 'd0;
    mem[13517] = 'd0;
    mem[13518] = 'd0;
    mem[13519] = 'd644;
    mem[13520] = 'd0;
    mem[13521] = 'd956;
    mem[13522] = 'd0;
    mem[13523] = 'd0;
    mem[13524] = 'd0;
    mem[13525] = 'd600;
    mem[13526] = 'd0;
    mem[13527] = 'd920;
    mem[13528] = 'd0;
    mem[13529] = 'd0;
    mem[13530] = 'd0;
    mem[13531] = 'd532;
    mem[13532] = 'd0;
    mem[13533] = 'd872;
    mem[13534] = 'd0;
    mem[13535] = 'd0;
    mem[13536] = 'd0;
    mem[13537] = 'd472;
    mem[13538] = 'd0;
    mem[13539] = 'd836;
    mem[13540] = 'd0;
    mem[13541] = 'd0;
    mem[13542] = 'd0;
    mem[13543] = 'd880;
    mem[13544] = 'd0;
    mem[13545] = 'd964;
    mem[13546] = 'd0;
    mem[13547] = 'd0;
    mem[13548] = 'd0;
    mem[13549] = 'd1020;
    mem[13550] = 'd0;
    mem[13551] = 'd1020;
    mem[13552] = 'd0;
    mem[13553] = 'd0;
    mem[13554] = 'd0;
    mem[13555] = 'd1020;
    mem[13556] = 'd0;
    mem[13557] = 'd1020;
    mem[13558] = 'd0;
    mem[13559] = 'd0;
    mem[13560] = 'd0;
    mem[13561] = 'd1020;
    mem[13562] = 'd0;
    mem[13563] = 'd1020;
    mem[13564] = 'd0;
    mem[13565] = 'd0;
    mem[13566] = 'd0;
    mem[13567] = 'd1020;
    mem[13568] = 'd0;
    mem[13569] = 'd1020;
    mem[13570] = 'd0;
    mem[13571] = 'd0;
    mem[13572] = 'd0;
    mem[13573] = 'd0;
    mem[13574] = 'd1020;
    mem[13575] = 'd0;
    mem[13576] = 'd1020;
    mem[13577] = 'd0;
    mem[13578] = 'd0;
    mem[13579] = 'd0;
    mem[13580] = 'd1020;
    mem[13581] = 'd0;
    mem[13582] = 'd1020;
    mem[13583] = 'd0;
    mem[13584] = 'd0;
    mem[13585] = 'd0;
    mem[13586] = 'd1020;
    mem[13587] = 'd0;
    mem[13588] = 'd1020;
    mem[13589] = 'd0;
    mem[13590] = 'd0;
    mem[13591] = 'd0;
    mem[13592] = 'd1016;
    mem[13593] = 'd0;
    mem[13594] = 'd1020;
    mem[13595] = 'd0;
    mem[13596] = 'd0;
    mem[13597] = 'd0;
    mem[13598] = 'd424;
    mem[13599] = 'd0;
    mem[13600] = 'd668;
    mem[13601] = 'd0;
    mem[13602] = 'd0;
    mem[13603] = 'd0;
    mem[13604] = 'd20;
    mem[13605] = 'd0;
    mem[13606] = 'd476;
    mem[13607] = 'd0;
    mem[13608] = 'd0;
    mem[13609] = 'd0;
    mem[13610] = 'd40;
    mem[13611] = 'd0;
    mem[13612] = 'd540;
    mem[13613] = 'd0;
    mem[13614] = 'd0;
    mem[13615] = 'd0;
    mem[13616] = 'd60;
    mem[13617] = 'd0;
    mem[13618] = 'd600;
    mem[13619] = 'd0;
    mem[13620] = 'd0;
    mem[13621] = 'd0;
    mem[13622] = 'd80;
    mem[13623] = 'd0;
    mem[13624] = 'd640;
    mem[13625] = 'd0;
    mem[13626] = 'd0;
    mem[13627] = 'd0;
    mem[13628] = 'd88;
    mem[13629] = 'd0;
    mem[13630] = 'd664;
    mem[13631] = 'd0;
    mem[13632] = 'd0;
    mem[13633] = 'd0;
    mem[13634] = 'd92;
    mem[13635] = 'd0;
    mem[13636] = 'd684;
    mem[13637] = 'd0;
    mem[13638] = 'd0;
    mem[13639] = 'd0;
    mem[13640] = 'd96;
    mem[13641] = 'd0;
    mem[13642] = 'd700;
    mem[13643] = 'd0;
    mem[13644] = 'd0;
    mem[13645] = 'd0;
    mem[13646] = 'd108;
    mem[13647] = 'd0;
    mem[13648] = 'd712;
    mem[13649] = 'd0;
    mem[13650] = 'd0;
    mem[13651] = 'd0;
    mem[13652] = 'd124;
    mem[13653] = 'd0;
    mem[13654] = 'd720;
    mem[13655] = 'd0;
    mem[13656] = 'd0;
    mem[13657] = 'd0;
    mem[13658] = 'd144;
    mem[13659] = 'd0;
    mem[13660] = 'd732;
    mem[13661] = 'd0;
    mem[13662] = 'd0;
    mem[13663] = 'd0;
    mem[13664] = 'd176;
    mem[13665] = 'd0;
    mem[13666] = 'd752;
    mem[13667] = 'd0;
    mem[13668] = 'd0;
    mem[13669] = 'd0;
    mem[13670] = 'd208;
    mem[13671] = 'd0;
    mem[13672] = 'd780;
    mem[13673] = 'd0;
    mem[13674] = 'd0;
    mem[13675] = 'd0;
    mem[13676] = 'd216;
    mem[13677] = 'd0;
    mem[13678] = 'd776;
    mem[13679] = 'd0;
    mem[13680] = 'd0;
    mem[13681] = 'd0;
    mem[13682] = 'd212;
    mem[13683] = 'd0;
    mem[13684] = 'd756;
    mem[13685] = 'd0;
    mem[13686] = 'd0;
    mem[13687] = 'd0;
    mem[13688] = 'd216;
    mem[13689] = 'd0;
    mem[13690] = 'd756;
    mem[13691] = 'd0;
    mem[13692] = 'd0;
    mem[13693] = 'd0;
    mem[13694] = 'd212;
    mem[13695] = 'd0;
    mem[13696] = 'd768;
    mem[13697] = 'd0;
    mem[13698] = 'd0;
    mem[13699] = 'd0;
    mem[13700] = 'd204;
    mem[13701] = 'd0;
    mem[13702] = 'd776;
    mem[13703] = 'd0;
    mem[13704] = 'd0;
    mem[13705] = 'd0;
    mem[13706] = 'd172;
    mem[13707] = 'd0;
    mem[13708] = 'd752;
    mem[13709] = 'd0;
    mem[13710] = 'd0;
    mem[13711] = 'd0;
    mem[13712] = 'd144;
    mem[13713] = 'd0;
    mem[13714] = 'd732;
    mem[13715] = 'd0;
    mem[13716] = 'd0;
    mem[13717] = 'd0;
    mem[13718] = 'd124;
    mem[13719] = 'd0;
    mem[13720] = 'd720;
    mem[13721] = 'd0;
    mem[13722] = 'd0;
    mem[13723] = 'd0;
    mem[13724] = 'd112;
    mem[13725] = 'd0;
    mem[13726] = 'd712;
    mem[13727] = 'd0;
    mem[13728] = 'd0;
    mem[13729] = 'd0;
    mem[13730] = 'd100;
    mem[13731] = 'd0;
    mem[13732] = 'd700;
    mem[13733] = 'd0;
    mem[13734] = 'd0;
    mem[13735] = 'd0;
    mem[13736] = 'd92;
    mem[13737] = 'd0;
    mem[13738] = 'd684;
    mem[13739] = 'd0;
    mem[13740] = 'd0;
    mem[13741] = 'd0;
    mem[13742] = 'd88;
    mem[13743] = 'd0;
    mem[13744] = 'd668;
    mem[13745] = 'd0;
    mem[13746] = 'd0;
    mem[13747] = 'd0;
    mem[13748] = 'd80;
    mem[13749] = 'd0;
    mem[13750] = 'd640;
    mem[13751] = 'd0;
    mem[13752] = 'd0;
    mem[13753] = 'd0;
    mem[13754] = 'd64;
    mem[13755] = 'd0;
    mem[13756] = 'd604;
    mem[13757] = 'd0;
    mem[13758] = 'd0;
    mem[13759] = 'd0;
    mem[13760] = 'd44;
    mem[13761] = 'd0;
    mem[13762] = 'd548;
    mem[13763] = 'd0;
    mem[13764] = 'd0;
    mem[13765] = 'd0;
    mem[13766] = 'd20;
    mem[13767] = 'd0;
    mem[13768] = 'd480;
    mem[13769] = 'd0;
    mem[13770] = 'd0;
    mem[13771] = 'd0;
    mem[13772] = 'd408;
    mem[13773] = 'd0;
    mem[13774] = 'd660;
    mem[13775] = 'd0;
    mem[13776] = 'd0;
    mem[13777] = 'd0;
    mem[13778] = 'd1016;
    mem[13779] = 'd0;
    mem[13780] = 'd1020;
    mem[13781] = 'd0;
    mem[13782] = 'd0;
    mem[13783] = 'd0;
    mem[13784] = 'd1020;
    mem[13785] = 'd0;
    mem[13786] = 'd1020;
    mem[13787] = 'd0;
    mem[13788] = 'd0;
    mem[13789] = 'd0;
    mem[13790] = 'd1020;
    mem[13791] = 'd0;
    mem[13792] = 'd1020;
    mem[13793] = 'd0;
    mem[13794] = 'd0;
    mem[13795] = 'd0;
    mem[13796] = 'd1020;
    mem[13797] = 'd0;
    mem[13798] = 'd1020;
    mem[13799] = 'd0;
    mem[13800] = 'd0;
    mem[13801] = 'd0;
    mem[13802] = 'd1020;
    mem[13803] = 'd0;
    mem[13804] = 'd1020;
    mem[13805] = 'd0;
    mem[13806] = 'd0;
    mem[13807] = 'd1020;
    mem[13808] = 'd0;
    mem[13809] = 'd1020;
    mem[13810] = 'd0;
    mem[13811] = 'd0;
    mem[13812] = 'd0;
    mem[13813] = 'd1020;
    mem[13814] = 'd0;
    mem[13815] = 'd1020;
    mem[13816] = 'd0;
    mem[13817] = 'd0;
    mem[13818] = 'd0;
    mem[13819] = 'd1020;
    mem[13820] = 'd0;
    mem[13821] = 'd1020;
    mem[13822] = 'd0;
    mem[13823] = 'd0;
    mem[13824] = 'd0;
    mem[13825] = 'd1020;
    mem[13826] = 'd0;
    mem[13827] = 'd1020;
    mem[13828] = 'd0;
    mem[13829] = 'd0;
    mem[13830] = 'd0;
    mem[13831] = 'd668;
    mem[13832] = 'd0;
    mem[13833] = 'd896;
    mem[13834] = 'd0;
    mem[13835] = 'd0;
    mem[13836] = 'd0;
    mem[13837] = 'd476;
    mem[13838] = 'd0;
    mem[13839] = 'd844;
    mem[13840] = 'd0;
    mem[13841] = 'd0;
    mem[13842] = 'd0;
    mem[13843] = 'd540;
    mem[13844] = 'd0;
    mem[13845] = 'd876;
    mem[13846] = 'd0;
    mem[13847] = 'd0;
    mem[13848] = 'd0;
    mem[13849] = 'd600;
    mem[13850] = 'd0;
    mem[13851] = 'd920;
    mem[13852] = 'd0;
    mem[13853] = 'd0;
    mem[13854] = 'd0;
    mem[13855] = 'd640;
    mem[13856] = 'd0;
    mem[13857] = 'd956;
    mem[13858] = 'd0;
    mem[13859] = 'd0;
    mem[13860] = 'd0;
    mem[13861] = 'd664;
    mem[13862] = 'd0;
    mem[13863] = 'd980;
    mem[13864] = 'd0;
    mem[13865] = 'd0;
    mem[13866] = 'd0;
    mem[13867] = 'd684;
    mem[13868] = 'd0;
    mem[13869] = 'd996;
    mem[13870] = 'd0;
    mem[13871] = 'd0;
    mem[13872] = 'd0;
    mem[13873] = 'd700;
    mem[13874] = 'd0;
    mem[13875] = 'd1012;
    mem[13876] = 'd0;
    mem[13877] = 'd0;
    mem[13878] = 'd0;
    mem[13879] = 'd712;
    mem[13880] = 'd0;
    mem[13881] = 'd1020;
    mem[13882] = 'd0;
    mem[13883] = 'd0;
    mem[13884] = 'd0;
    mem[13885] = 'd720;
    mem[13886] = 'd0;
    mem[13887] = 'd1020;
    mem[13888] = 'd0;
    mem[13889] = 'd0;
    mem[13890] = 'd0;
    mem[13891] = 'd732;
    mem[13892] = 'd0;
    mem[13893] = 'd1020;
    mem[13894] = 'd0;
    mem[13895] = 'd0;
    mem[13896] = 'd0;
    mem[13897] = 'd752;
    mem[13898] = 'd0;
    mem[13899] = 'd1020;
    mem[13900] = 'd0;
    mem[13901] = 'd0;
    mem[13902] = 'd0;
    mem[13903] = 'd780;
    mem[13904] = 'd0;
    mem[13905] = 'd1012;
    mem[13906] = 'd0;
    mem[13907] = 'd0;
    mem[13908] = 'd0;
    mem[13909] = 'd776;
    mem[13910] = 'd0;
    mem[13911] = 'd984;
    mem[13912] = 'd0;
    mem[13913] = 'd0;
    mem[13914] = 'd0;
    mem[13915] = 'd756;
    mem[13916] = 'd0;
    mem[13917] = 'd960;
    mem[13918] = 'd0;
    mem[13919] = 'd0;
    mem[13920] = 'd0;
    mem[13921] = 'd756;
    mem[13922] = 'd0;
    mem[13923] = 'd960;
    mem[13924] = 'd0;
    mem[13925] = 'd0;
    mem[13926] = 'd0;
    mem[13927] = 'd768;
    mem[13928] = 'd0;
    mem[13929] = 'd976;
    mem[13930] = 'd0;
    mem[13931] = 'd0;
    mem[13932] = 'd0;
    mem[13933] = 'd776;
    mem[13934] = 'd0;
    mem[13935] = 'd1012;
    mem[13936] = 'd0;
    mem[13937] = 'd0;
    mem[13938] = 'd0;
    mem[13939] = 'd752;
    mem[13940] = 'd0;
    mem[13941] = 'd1020;
    mem[13942] = 'd0;
    mem[13943] = 'd0;
    mem[13944] = 'd0;
    mem[13945] = 'd732;
    mem[13946] = 'd0;
    mem[13947] = 'd1020;
    mem[13948] = 'd0;
    mem[13949] = 'd0;
    mem[13950] = 'd0;
    mem[13951] = 'd720;
    mem[13952] = 'd0;
    mem[13953] = 'd1020;
    mem[13954] = 'd0;
    mem[13955] = 'd0;
    mem[13956] = 'd0;
    mem[13957] = 'd712;
    mem[13958] = 'd0;
    mem[13959] = 'd1020;
    mem[13960] = 'd0;
    mem[13961] = 'd0;
    mem[13962] = 'd0;
    mem[13963] = 'd700;
    mem[13964] = 'd0;
    mem[13965] = 'd1012;
    mem[13966] = 'd0;
    mem[13967] = 'd0;
    mem[13968] = 'd0;
    mem[13969] = 'd684;
    mem[13970] = 'd0;
    mem[13971] = 'd1000;
    mem[13972] = 'd0;
    mem[13973] = 'd0;
    mem[13974] = 'd0;
    mem[13975] = 'd668;
    mem[13976] = 'd0;
    mem[13977] = 'd984;
    mem[13978] = 'd0;
    mem[13979] = 'd0;
    mem[13980] = 'd0;
    mem[13981] = 'd640;
    mem[13982] = 'd0;
    mem[13983] = 'd956;
    mem[13984] = 'd0;
    mem[13985] = 'd0;
    mem[13986] = 'd0;
    mem[13987] = 'd604;
    mem[13988] = 'd0;
    mem[13989] = 'd924;
    mem[13990] = 'd0;
    mem[13991] = 'd0;
    mem[13992] = 'd0;
    mem[13993] = 'd548;
    mem[13994] = 'd0;
    mem[13995] = 'd880;
    mem[13996] = 'd0;
    mem[13997] = 'd0;
    mem[13998] = 'd0;
    mem[13999] = 'd480;
    mem[14000] = 'd0;
    mem[14001] = 'd844;
    mem[14002] = 'd0;
    mem[14003] = 'd0;
    mem[14004] = 'd0;
    mem[14005] = 'd660;
    mem[14006] = 'd0;
    mem[14007] = 'd892;
    mem[14008] = 'd0;
    mem[14009] = 'd0;
    mem[14010] = 'd0;
    mem[14011] = 'd1020;
    mem[14012] = 'd0;
    mem[14013] = 'd1020;
    mem[14014] = 'd0;
    mem[14015] = 'd0;
    mem[14016] = 'd0;
    mem[14017] = 'd1020;
    mem[14018] = 'd0;
    mem[14019] = 'd1020;
    mem[14020] = 'd0;
    mem[14021] = 'd0;
    mem[14022] = 'd0;
    mem[14023] = 'd1020;
    mem[14024] = 'd0;
    mem[14025] = 'd1020;
    mem[14026] = 'd0;
    mem[14027] = 'd0;
    mem[14028] = 'd0;
    mem[14029] = 'd1020;
    mem[14030] = 'd0;
    mem[14031] = 'd1020;
    mem[14032] = 'd0;
    mem[14033] = 'd0;
    mem[14034] = 'd0;
    mem[14035] = 'd1020;
    mem[14036] = 'd0;
    mem[14037] = 'd1020;
    mem[14038] = 'd0;
    mem[14039] = 'd0;
    mem[14040] = 'd0;
    mem[14041] = 'd0;
    mem[14042] = 'd1020;
    mem[14043] = 'd0;
    mem[14044] = 'd1020;
    mem[14045] = 'd0;
    mem[14046] = 'd0;
    mem[14047] = 'd0;
    mem[14048] = 'd1020;
    mem[14049] = 'd0;
    mem[14050] = 'd1020;
    mem[14051] = 'd0;
    mem[14052] = 'd0;
    mem[14053] = 'd0;
    mem[14054] = 'd1020;
    mem[14055] = 'd0;
    mem[14056] = 'd1020;
    mem[14057] = 'd0;
    mem[14058] = 'd0;
    mem[14059] = 'd0;
    mem[14060] = 'd1016;
    mem[14061] = 'd0;
    mem[14062] = 'd1020;
    mem[14063] = 'd0;
    mem[14064] = 'd0;
    mem[14065] = 'd0;
    mem[14066] = 'd948;
    mem[14067] = 'd0;
    mem[14068] = 'd976;
    mem[14069] = 'd0;
    mem[14070] = 'd0;
    mem[14071] = 'd0;
    mem[14072] = 'd220;
    mem[14073] = 'd0;
    mem[14074] = 'd540;
    mem[14075] = 'd0;
    mem[14076] = 'd0;
    mem[14077] = 'd0;
    mem[14078] = 'd24;
    mem[14079] = 'd0;
    mem[14080] = 'd488;
    mem[14081] = 'd0;
    mem[14082] = 'd0;
    mem[14083] = 'd0;
    mem[14084] = 'd44;
    mem[14085] = 'd0;
    mem[14086] = 'd548;
    mem[14087] = 'd0;
    mem[14088] = 'd0;
    mem[14089] = 'd0;
    mem[14090] = 'd60;
    mem[14091] = 'd0;
    mem[14092] = 'd596;
    mem[14093] = 'd0;
    mem[14094] = 'd0;
    mem[14095] = 'd0;
    mem[14096] = 'd76;
    mem[14097] = 'd0;
    mem[14098] = 'd632;
    mem[14099] = 'd0;
    mem[14100] = 'd0;
    mem[14101] = 'd0;
    mem[14102] = 'd84;
    mem[14103] = 'd0;
    mem[14104] = 'd656;
    mem[14105] = 'd0;
    mem[14106] = 'd0;
    mem[14107] = 'd0;
    mem[14108] = 'd88;
    mem[14109] = 'd0;
    mem[14110] = 'd672;
    mem[14111] = 'd0;
    mem[14112] = 'd0;
    mem[14113] = 'd0;
    mem[14114] = 'd92;
    mem[14115] = 'd0;
    mem[14116] = 'd688;
    mem[14117] = 'd0;
    mem[14118] = 'd0;
    mem[14119] = 'd0;
    mem[14120] = 'd96;
    mem[14121] = 'd0;
    mem[14122] = 'd696;
    mem[14123] = 'd0;
    mem[14124] = 'd0;
    mem[14125] = 'd0;
    mem[14126] = 'd104;
    mem[14127] = 'd0;
    mem[14128] = 'd704;
    mem[14129] = 'd0;
    mem[14130] = 'd0;
    mem[14131] = 'd0;
    mem[14132] = 'd116;
    mem[14133] = 'd0;
    mem[14134] = 'd712;
    mem[14135] = 'd0;
    mem[14136] = 'd0;
    mem[14137] = 'd0;
    mem[14138] = 'd128;
    mem[14139] = 'd0;
    mem[14140] = 'd716;
    mem[14141] = 'd0;
    mem[14142] = 'd0;
    mem[14143] = 'd0;
    mem[14144] = 'd132;
    mem[14145] = 'd0;
    mem[14146] = 'd716;
    mem[14147] = 'd0;
    mem[14148] = 'd0;
    mem[14149] = 'd0;
    mem[14150] = 'd132;
    mem[14151] = 'd0;
    mem[14152] = 'd720;
    mem[14153] = 'd0;
    mem[14154] = 'd0;
    mem[14155] = 'd0;
    mem[14156] = 'd132;
    mem[14157] = 'd0;
    mem[14158] = 'd716;
    mem[14159] = 'd0;
    mem[14160] = 'd0;
    mem[14161] = 'd0;
    mem[14162] = 'd132;
    mem[14163] = 'd0;
    mem[14164] = 'd716;
    mem[14165] = 'd0;
    mem[14166] = 'd0;
    mem[14167] = 'd0;
    mem[14168] = 'd128;
    mem[14169] = 'd0;
    mem[14170] = 'd716;
    mem[14171] = 'd0;
    mem[14172] = 'd0;
    mem[14173] = 'd0;
    mem[14174] = 'd120;
    mem[14175] = 'd0;
    mem[14176] = 'd712;
    mem[14177] = 'd0;
    mem[14178] = 'd0;
    mem[14179] = 'd0;
    mem[14180] = 'd104;
    mem[14181] = 'd0;
    mem[14182] = 'd704;
    mem[14183] = 'd0;
    mem[14184] = 'd0;
    mem[14185] = 'd0;
    mem[14186] = 'd92;
    mem[14187] = 'd0;
    mem[14188] = 'd696;
    mem[14189] = 'd0;
    mem[14190] = 'd0;
    mem[14191] = 'd0;
    mem[14192] = 'd92;
    mem[14193] = 'd0;
    mem[14194] = 'd688;
    mem[14195] = 'd0;
    mem[14196] = 'd0;
    mem[14197] = 'd0;
    mem[14198] = 'd88;
    mem[14199] = 'd0;
    mem[14200] = 'd676;
    mem[14201] = 'd0;
    mem[14202] = 'd0;
    mem[14203] = 'd0;
    mem[14204] = 'd88;
    mem[14205] = 'd0;
    mem[14206] = 'd660;
    mem[14207] = 'd0;
    mem[14208] = 'd0;
    mem[14209] = 'd0;
    mem[14210] = 'd80;
    mem[14211] = 'd0;
    mem[14212] = 'd636;
    mem[14213] = 'd0;
    mem[14214] = 'd0;
    mem[14215] = 'd0;
    mem[14216] = 'd68;
    mem[14217] = 'd0;
    mem[14218] = 'd600;
    mem[14219] = 'd0;
    mem[14220] = 'd0;
    mem[14221] = 'd0;
    mem[14222] = 'd48;
    mem[14223] = 'd0;
    mem[14224] = 'd552;
    mem[14225] = 'd0;
    mem[14226] = 'd0;
    mem[14227] = 'd0;
    mem[14228] = 'd24;
    mem[14229] = 'd0;
    mem[14230] = 'd492;
    mem[14231] = 'd0;
    mem[14232] = 'd0;
    mem[14233] = 'd0;
    mem[14234] = 'd192;
    mem[14235] = 'd0;
    mem[14236] = 'd520;
    mem[14237] = 'd0;
    mem[14238] = 'd0;
    mem[14239] = 'd0;
    mem[14240] = 'd936;
    mem[14241] = 'd0;
    mem[14242] = 'd964;
    mem[14243] = 'd0;
    mem[14244] = 'd0;
    mem[14245] = 'd0;
    mem[14246] = 'd1016;
    mem[14247] = 'd0;
    mem[14248] = 'd1020;
    mem[14249] = 'd0;
    mem[14250] = 'd0;
    mem[14251] = 'd0;
    mem[14252] = 'd1020;
    mem[14253] = 'd0;
    mem[14254] = 'd1020;
    mem[14255] = 'd0;
    mem[14256] = 'd0;
    mem[14257] = 'd0;
    mem[14258] = 'd1020;
    mem[14259] = 'd0;
    mem[14260] = 'd1020;
    mem[14261] = 'd0;
    mem[14262] = 'd0;
    mem[14263] = 'd0;
    mem[14264] = 'd1020;
    mem[14265] = 'd0;
    mem[14266] = 'd1020;
    mem[14267] = 'd0;
    mem[14268] = 'd0;
    mem[14269] = 'd0;
    mem[14270] = 'd1020;
    mem[14271] = 'd0;
    mem[14272] = 'd1020;
    mem[14273] = 'd0;
    mem[14274] = 'd0;
    mem[14275] = 'd1020;
    mem[14276] = 'd0;
    mem[14277] = 'd1020;
    mem[14278] = 'd0;
    mem[14279] = 'd0;
    mem[14280] = 'd0;
    mem[14281] = 'd1020;
    mem[14282] = 'd0;
    mem[14283] = 'd1020;
    mem[14284] = 'd0;
    mem[14285] = 'd0;
    mem[14286] = 'd0;
    mem[14287] = 'd1020;
    mem[14288] = 'd0;
    mem[14289] = 'd1020;
    mem[14290] = 'd0;
    mem[14291] = 'd0;
    mem[14292] = 'd0;
    mem[14293] = 'd1020;
    mem[14294] = 'd0;
    mem[14295] = 'd1020;
    mem[14296] = 'd0;
    mem[14297] = 'd0;
    mem[14298] = 'd0;
    mem[14299] = 'd976;
    mem[14300] = 'd0;
    mem[14301] = 'd1000;
    mem[14302] = 'd0;
    mem[14303] = 'd0;
    mem[14304] = 'd0;
    mem[14305] = 'd540;
    mem[14306] = 'd0;
    mem[14307] = 'd844;
    mem[14308] = 'd0;
    mem[14309] = 'd0;
    mem[14310] = 'd0;
    mem[14311] = 'd488;
    mem[14312] = 'd0;
    mem[14313] = 'd848;
    mem[14314] = 'd0;
    mem[14315] = 'd0;
    mem[14316] = 'd0;
    mem[14317] = 'd548;
    mem[14318] = 'd0;
    mem[14319] = 'd880;
    mem[14320] = 'd0;
    mem[14321] = 'd0;
    mem[14322] = 'd0;
    mem[14323] = 'd596;
    mem[14324] = 'd0;
    mem[14325] = 'd916;
    mem[14326] = 'd0;
    mem[14327] = 'd0;
    mem[14328] = 'd0;
    mem[14329] = 'd632;
    mem[14330] = 'd0;
    mem[14331] = 'd952;
    mem[14332] = 'd0;
    mem[14333] = 'd0;
    mem[14334] = 'd0;
    mem[14335] = 'd656;
    mem[14336] = 'd0;
    mem[14337] = 'd972;
    mem[14338] = 'd0;
    mem[14339] = 'd0;
    mem[14340] = 'd0;
    mem[14341] = 'd672;
    mem[14342] = 'd0;
    mem[14343] = 'd992;
    mem[14344] = 'd0;
    mem[14345] = 'd0;
    mem[14346] = 'd0;
    mem[14347] = 'd688;
    mem[14348] = 'd0;
    mem[14349] = 'd1004;
    mem[14350] = 'd0;
    mem[14351] = 'd0;
    mem[14352] = 'd0;
    mem[14353] = 'd696;
    mem[14354] = 'd0;
    mem[14355] = 'd1016;
    mem[14356] = 'd0;
    mem[14357] = 'd0;
    mem[14358] = 'd0;
    mem[14359] = 'd704;
    mem[14360] = 'd0;
    mem[14361] = 'd1020;
    mem[14362] = 'd0;
    mem[14363] = 'd0;
    mem[14364] = 'd0;
    mem[14365] = 'd712;
    mem[14366] = 'd0;
    mem[14367] = 'd1020;
    mem[14368] = 'd0;
    mem[14369] = 'd0;
    mem[14370] = 'd0;
    mem[14371] = 'd716;
    mem[14372] = 'd0;
    mem[14373] = 'd1020;
    mem[14374] = 'd0;
    mem[14375] = 'd0;
    mem[14376] = 'd0;
    mem[14377] = 'd716;
    mem[14378] = 'd0;
    mem[14379] = 'd1020;
    mem[14380] = 'd0;
    mem[14381] = 'd0;
    mem[14382] = 'd0;
    mem[14383] = 'd720;
    mem[14384] = 'd0;
    mem[14385] = 'd1020;
    mem[14386] = 'd0;
    mem[14387] = 'd0;
    mem[14388] = 'd0;
    mem[14389] = 'd716;
    mem[14390] = 'd0;
    mem[14391] = 'd1020;
    mem[14392] = 'd0;
    mem[14393] = 'd0;
    mem[14394] = 'd0;
    mem[14395] = 'd716;
    mem[14396] = 'd0;
    mem[14397] = 'd1020;
    mem[14398] = 'd0;
    mem[14399] = 'd0;
    mem[14400] = 'd0;
    mem[14401] = 'd716;
    mem[14402] = 'd0;
    mem[14403] = 'd1020;
    mem[14404] = 'd0;
    mem[14405] = 'd0;
    mem[14406] = 'd0;
    mem[14407] = 'd712;
    mem[14408] = 'd0;
    mem[14409] = 'd1020;
    mem[14410] = 'd0;
    mem[14411] = 'd0;
    mem[14412] = 'd0;
    mem[14413] = 'd704;
    mem[14414] = 'd0;
    mem[14415] = 'd1020;
    mem[14416] = 'd0;
    mem[14417] = 'd0;
    mem[14418] = 'd0;
    mem[14419] = 'd696;
    mem[14420] = 'd0;
    mem[14421] = 'd1016;
    mem[14422] = 'd0;
    mem[14423] = 'd0;
    mem[14424] = 'd0;
    mem[14425] = 'd688;
    mem[14426] = 'd0;
    mem[14427] = 'd1008;
    mem[14428] = 'd0;
    mem[14429] = 'd0;
    mem[14430] = 'd0;
    mem[14431] = 'd676;
    mem[14432] = 'd0;
    mem[14433] = 'd992;
    mem[14434] = 'd0;
    mem[14435] = 'd0;
    mem[14436] = 'd0;
    mem[14437] = 'd660;
    mem[14438] = 'd0;
    mem[14439] = 'd976;
    mem[14440] = 'd0;
    mem[14441] = 'd0;
    mem[14442] = 'd0;
    mem[14443] = 'd636;
    mem[14444] = 'd0;
    mem[14445] = 'd952;
    mem[14446] = 'd0;
    mem[14447] = 'd0;
    mem[14448] = 'd0;
    mem[14449] = 'd600;
    mem[14450] = 'd0;
    mem[14451] = 'd920;
    mem[14452] = 'd0;
    mem[14453] = 'd0;
    mem[14454] = 'd0;
    mem[14455] = 'd552;
    mem[14456] = 'd0;
    mem[14457] = 'd884;
    mem[14458] = 'd0;
    mem[14459] = 'd0;
    mem[14460] = 'd0;
    mem[14461] = 'd492;
    mem[14462] = 'd0;
    mem[14463] = 'd852;
    mem[14464] = 'd0;
    mem[14465] = 'd0;
    mem[14466] = 'd0;
    mem[14467] = 'd520;
    mem[14468] = 'd0;
    mem[14469] = 'd836;
    mem[14470] = 'd0;
    mem[14471] = 'd0;
    mem[14472] = 'd0;
    mem[14473] = 'd964;
    mem[14474] = 'd0;
    mem[14475] = 'd996;
    mem[14476] = 'd0;
    mem[14477] = 'd0;
    mem[14478] = 'd0;
    mem[14479] = 'd1020;
    mem[14480] = 'd0;
    mem[14481] = 'd1020;
    mem[14482] = 'd0;
    mem[14483] = 'd0;
    mem[14484] = 'd0;
    mem[14485] = 'd1020;
    mem[14486] = 'd0;
    mem[14487] = 'd1020;
    mem[14488] = 'd0;
    mem[14489] = 'd0;
    mem[14490] = 'd0;
    mem[14491] = 'd1020;
    mem[14492] = 'd0;
    mem[14493] = 'd1020;
    mem[14494] = 'd0;
    mem[14495] = 'd0;
    mem[14496] = 'd0;
    mem[14497] = 'd1020;
    mem[14498] = 'd0;
    mem[14499] = 'd1020;
    mem[14500] = 'd0;
    mem[14501] = 'd0;
    mem[14502] = 'd0;
    mem[14503] = 'd1020;
    mem[14504] = 'd0;
    mem[14505] = 'd1020;
    mem[14506] = 'd0;
    mem[14507] = 'd0;
    mem[14508] = 'd0;
    mem[14509] = 'd0;
    mem[14510] = 'd1020;
    mem[14511] = 'd0;
    mem[14512] = 'd1020;
    mem[14513] = 'd0;
    mem[14514] = 'd0;
    mem[14515] = 'd0;
    mem[14516] = 'd1020;
    mem[14517] = 'd0;
    mem[14518] = 'd1020;
    mem[14519] = 'd0;
    mem[14520] = 'd0;
    mem[14521] = 'd0;
    mem[14522] = 'd1020;
    mem[14523] = 'd0;
    mem[14524] = 'd1020;
    mem[14525] = 'd0;
    mem[14526] = 'd0;
    mem[14527] = 'd0;
    mem[14528] = 'd1020;
    mem[14529] = 'd0;
    mem[14530] = 'd1020;
    mem[14531] = 'd0;
    mem[14532] = 'd0;
    mem[14533] = 'd0;
    mem[14534] = 'd1016;
    mem[14535] = 'd0;
    mem[14536] = 'd1020;
    mem[14537] = 'd0;
    mem[14538] = 'd0;
    mem[14539] = 'd0;
    mem[14540] = 'd900;
    mem[14541] = 'd0;
    mem[14542] = 'd944;
    mem[14543] = 'd0;
    mem[14544] = 'd0;
    mem[14545] = 'd0;
    mem[14546] = 'd168;
    mem[14547] = 'd0;
    mem[14548] = 'd504;
    mem[14549] = 'd0;
    mem[14550] = 'd0;
    mem[14551] = 'd0;
    mem[14552] = 'd24;
    mem[14553] = 'd0;
    mem[14554] = 'd488;
    mem[14555] = 'd0;
    mem[14556] = 'd0;
    mem[14557] = 'd0;
    mem[14558] = 'd40;
    mem[14559] = 'd0;
    mem[14560] = 'd540;
    mem[14561] = 'd0;
    mem[14562] = 'd0;
    mem[14563] = 'd0;
    mem[14564] = 'd56;
    mem[14565] = 'd0;
    mem[14566] = 'd584;
    mem[14567] = 'd0;
    mem[14568] = 'd0;
    mem[14569] = 'd0;
    mem[14570] = 'd72;
    mem[14571] = 'd0;
    mem[14572] = 'd620;
    mem[14573] = 'd0;
    mem[14574] = 'd0;
    mem[14575] = 'd0;
    mem[14576] = 'd80;
    mem[14577] = 'd0;
    mem[14578] = 'd644;
    mem[14579] = 'd0;
    mem[14580] = 'd0;
    mem[14581] = 'd0;
    mem[14582] = 'd88;
    mem[14583] = 'd0;
    mem[14584] = 'd660;
    mem[14585] = 'd0;
    mem[14586] = 'd0;
    mem[14587] = 'd0;
    mem[14588] = 'd88;
    mem[14589] = 'd0;
    mem[14590] = 'd672;
    mem[14591] = 'd0;
    mem[14592] = 'd0;
    mem[14593] = 'd0;
    mem[14594] = 'd92;
    mem[14595] = 'd0;
    mem[14596] = 'd680;
    mem[14597] = 'd0;
    mem[14598] = 'd0;
    mem[14599] = 'd0;
    mem[14600] = 'd92;
    mem[14601] = 'd0;
    mem[14602] = 'd688;
    mem[14603] = 'd0;
    mem[14604] = 'd0;
    mem[14605] = 'd0;
    mem[14606] = 'd92;
    mem[14607] = 'd0;
    mem[14608] = 'd692;
    mem[14609] = 'd0;
    mem[14610] = 'd0;
    mem[14611] = 'd0;
    mem[14612] = 'd96;
    mem[14613] = 'd0;
    mem[14614] = 'd692;
    mem[14615] = 'd0;
    mem[14616] = 'd0;
    mem[14617] = 'd0;
    mem[14618] = 'd96;
    mem[14619] = 'd0;
    mem[14620] = 'd692;
    mem[14621] = 'd0;
    mem[14622] = 'd0;
    mem[14623] = 'd0;
    mem[14624] = 'd100;
    mem[14625] = 'd0;
    mem[14626] = 'd696;
    mem[14627] = 'd0;
    mem[14628] = 'd0;
    mem[14629] = 'd0;
    mem[14630] = 'd96;
    mem[14631] = 'd0;
    mem[14632] = 'd692;
    mem[14633] = 'd0;
    mem[14634] = 'd0;
    mem[14635] = 'd0;
    mem[14636] = 'd92;
    mem[14637] = 'd0;
    mem[14638] = 'd692;
    mem[14639] = 'd0;
    mem[14640] = 'd0;
    mem[14641] = 'd0;
    mem[14642] = 'd92;
    mem[14643] = 'd0;
    mem[14644] = 'd684;
    mem[14645] = 'd0;
    mem[14646] = 'd0;
    mem[14647] = 'd0;
    mem[14648] = 'd92;
    mem[14649] = 'd0;
    mem[14650] = 'd680;
    mem[14651] = 'd0;
    mem[14652] = 'd0;
    mem[14653] = 'd0;
    mem[14654] = 'd88;
    mem[14655] = 'd0;
    mem[14656] = 'd676;
    mem[14657] = 'd0;
    mem[14658] = 'd0;
    mem[14659] = 'd0;
    mem[14660] = 'd88;
    mem[14661] = 'd0;
    mem[14662] = 'd664;
    mem[14663] = 'd0;
    mem[14664] = 'd0;
    mem[14665] = 'd0;
    mem[14666] = 'd84;
    mem[14667] = 'd0;
    mem[14668] = 'd648;
    mem[14669] = 'd0;
    mem[14670] = 'd0;
    mem[14671] = 'd0;
    mem[14672] = 'd76;
    mem[14673] = 'd0;
    mem[14674] = 'd624;
    mem[14675] = 'd0;
    mem[14676] = 'd0;
    mem[14677] = 'd0;
    mem[14678] = 'd60;
    mem[14679] = 'd0;
    mem[14680] = 'd588;
    mem[14681] = 'd0;
    mem[14682] = 'd0;
    mem[14683] = 'd0;
    mem[14684] = 'd44;
    mem[14685] = 'd0;
    mem[14686] = 'd548;
    mem[14687] = 'd0;
    mem[14688] = 'd0;
    mem[14689] = 'd0;
    mem[14690] = 'd24;
    mem[14691] = 'd0;
    mem[14692] = 'd492;
    mem[14693] = 'd0;
    mem[14694] = 'd0;
    mem[14695] = 'd0;
    mem[14696] = 'd144;
    mem[14697] = 'd0;
    mem[14698] = 'd496;
    mem[14699] = 'd0;
    mem[14700] = 'd0;
    mem[14701] = 'd0;
    mem[14702] = 'd892;
    mem[14703] = 'd0;
    mem[14704] = 'd940;
    mem[14705] = 'd0;
    mem[14706] = 'd0;
    mem[14707] = 'd0;
    mem[14708] = 'd1016;
    mem[14709] = 'd0;
    mem[14710] = 'd1020;
    mem[14711] = 'd0;
    mem[14712] = 'd0;
    mem[14713] = 'd0;
    mem[14714] = 'd1020;
    mem[14715] = 'd0;
    mem[14716] = 'd1020;
    mem[14717] = 'd0;
    mem[14718] = 'd0;
    mem[14719] = 'd0;
    mem[14720] = 'd1020;
    mem[14721] = 'd0;
    mem[14722] = 'd1020;
    mem[14723] = 'd0;
    mem[14724] = 'd0;
    mem[14725] = 'd0;
    mem[14726] = 'd1020;
    mem[14727] = 'd0;
    mem[14728] = 'd1020;
    mem[14729] = 'd0;
    mem[14730] = 'd0;
    mem[14731] = 'd0;
    mem[14732] = 'd1020;
    mem[14733] = 'd0;
    mem[14734] = 'd1020;
    mem[14735] = 'd0;
    mem[14736] = 'd0;
    mem[14737] = 'd0;
    mem[14738] = 'd1020;
    mem[14739] = 'd0;
    mem[14740] = 'd1020;
    mem[14741] = 'd0;
    mem[14742] = 'd0;
    mem[14743] = 'd1020;
    mem[14744] = 'd0;
    mem[14745] = 'd1020;
    mem[14746] = 'd0;
    mem[14747] = 'd0;
    mem[14748] = 'd0;
    mem[14749] = 'd1020;
    mem[14750] = 'd0;
    mem[14751] = 'd1020;
    mem[14752] = 'd0;
    mem[14753] = 'd0;
    mem[14754] = 'd0;
    mem[14755] = 'd1020;
    mem[14756] = 'd0;
    mem[14757] = 'd1020;
    mem[14758] = 'd0;
    mem[14759] = 'd0;
    mem[14760] = 'd0;
    mem[14761] = 'd1020;
    mem[14762] = 'd0;
    mem[14763] = 'd1020;
    mem[14764] = 'd0;
    mem[14765] = 'd0;
    mem[14766] = 'd0;
    mem[14767] = 'd1020;
    mem[14768] = 'd0;
    mem[14769] = 'd1020;
    mem[14770] = 'd0;
    mem[14771] = 'd0;
    mem[14772] = 'd0;
    mem[14773] = 'd944;
    mem[14774] = 'd0;
    mem[14775] = 'd988;
    mem[14776] = 'd0;
    mem[14777] = 'd0;
    mem[14778] = 'd0;
    mem[14779] = 'd504;
    mem[14780] = 'd0;
    mem[14781] = 'd824;
    mem[14782] = 'd0;
    mem[14783] = 'd0;
    mem[14784] = 'd0;
    mem[14785] = 'd488;
    mem[14786] = 'd0;
    mem[14787] = 'd852;
    mem[14788] = 'd0;
    mem[14789] = 'd0;
    mem[14790] = 'd0;
    mem[14791] = 'd540;
    mem[14792] = 'd0;
    mem[14793] = 'd880;
    mem[14794] = 'd0;
    mem[14795] = 'd0;
    mem[14796] = 'd0;
    mem[14797] = 'd584;
    mem[14798] = 'd0;
    mem[14799] = 'd908;
    mem[14800] = 'd0;
    mem[14801] = 'd0;
    mem[14802] = 'd0;
    mem[14803] = 'd620;
    mem[14804] = 'd0;
    mem[14805] = 'd940;
    mem[14806] = 'd0;
    mem[14807] = 'd0;
    mem[14808] = 'd0;
    mem[14809] = 'd644;
    mem[14810] = 'd0;
    mem[14811] = 'd960;
    mem[14812] = 'd0;
    mem[14813] = 'd0;
    mem[14814] = 'd0;
    mem[14815] = 'd660;
    mem[14816] = 'd0;
    mem[14817] = 'd980;
    mem[14818] = 'd0;
    mem[14819] = 'd0;
    mem[14820] = 'd0;
    mem[14821] = 'd672;
    mem[14822] = 'd0;
    mem[14823] = 'd996;
    mem[14824] = 'd0;
    mem[14825] = 'd0;
    mem[14826] = 'd0;
    mem[14827] = 'd680;
    mem[14828] = 'd0;
    mem[14829] = 'd1004;
    mem[14830] = 'd0;
    mem[14831] = 'd0;
    mem[14832] = 'd0;
    mem[14833] = 'd688;
    mem[14834] = 'd0;
    mem[14835] = 'd1012;
    mem[14836] = 'd0;
    mem[14837] = 'd0;
    mem[14838] = 'd0;
    mem[14839] = 'd692;
    mem[14840] = 'd0;
    mem[14841] = 'd1016;
    mem[14842] = 'd0;
    mem[14843] = 'd0;
    mem[14844] = 'd0;
    mem[14845] = 'd692;
    mem[14846] = 'd0;
    mem[14847] = 'd1016;
    mem[14848] = 'd0;
    mem[14849] = 'd0;
    mem[14850] = 'd0;
    mem[14851] = 'd692;
    mem[14852] = 'd0;
    mem[14853] = 'd1016;
    mem[14854] = 'd0;
    mem[14855] = 'd0;
    mem[14856] = 'd0;
    mem[14857] = 'd696;
    mem[14858] = 'd0;
    mem[14859] = 'd1016;
    mem[14860] = 'd0;
    mem[14861] = 'd0;
    mem[14862] = 'd0;
    mem[14863] = 'd692;
    mem[14864] = 'd0;
    mem[14865] = 'd1016;
    mem[14866] = 'd0;
    mem[14867] = 'd0;
    mem[14868] = 'd0;
    mem[14869] = 'd692;
    mem[14870] = 'd0;
    mem[14871] = 'd1016;
    mem[14872] = 'd0;
    mem[14873] = 'd0;
    mem[14874] = 'd0;
    mem[14875] = 'd684;
    mem[14876] = 'd0;
    mem[14877] = 'd1012;
    mem[14878] = 'd0;
    mem[14879] = 'd0;
    mem[14880] = 'd0;
    mem[14881] = 'd680;
    mem[14882] = 'd0;
    mem[14883] = 'd1004;
    mem[14884] = 'd0;
    mem[14885] = 'd0;
    mem[14886] = 'd0;
    mem[14887] = 'd676;
    mem[14888] = 'd0;
    mem[14889] = 'd996;
    mem[14890] = 'd0;
    mem[14891] = 'd0;
    mem[14892] = 'd0;
    mem[14893] = 'd664;
    mem[14894] = 'd0;
    mem[14895] = 'd984;
    mem[14896] = 'd0;
    mem[14897] = 'd0;
    mem[14898] = 'd0;
    mem[14899] = 'd648;
    mem[14900] = 'd0;
    mem[14901] = 'd968;
    mem[14902] = 'd0;
    mem[14903] = 'd0;
    mem[14904] = 'd0;
    mem[14905] = 'd624;
    mem[14906] = 'd0;
    mem[14907] = 'd940;
    mem[14908] = 'd0;
    mem[14909] = 'd0;
    mem[14910] = 'd0;
    mem[14911] = 'd588;
    mem[14912] = 'd0;
    mem[14913] = 'd912;
    mem[14914] = 'd0;
    mem[14915] = 'd0;
    mem[14916] = 'd0;
    mem[14917] = 'd548;
    mem[14918] = 'd0;
    mem[14919] = 'd884;
    mem[14920] = 'd0;
    mem[14921] = 'd0;
    mem[14922] = 'd0;
    mem[14923] = 'd492;
    mem[14924] = 'd0;
    mem[14925] = 'd852;
    mem[14926] = 'd0;
    mem[14927] = 'd0;
    mem[14928] = 'd0;
    mem[14929] = 'd496;
    mem[14930] = 'd0;
    mem[14931] = 'd828;
    mem[14932] = 'd0;
    mem[14933] = 'd0;
    mem[14934] = 'd0;
    mem[14935] = 'd940;
    mem[14936] = 'd0;
    mem[14937] = 'd988;
    mem[14938] = 'd0;
    mem[14939] = 'd0;
    mem[14940] = 'd0;
    mem[14941] = 'd1020;
    mem[14942] = 'd0;
    mem[14943] = 'd1020;
    mem[14944] = 'd0;
    mem[14945] = 'd0;
    mem[14946] = 'd0;
    mem[14947] = 'd1020;
    mem[14948] = 'd0;
    mem[14949] = 'd1020;
    mem[14950] = 'd0;
    mem[14951] = 'd0;
    mem[14952] = 'd0;
    mem[14953] = 'd1020;
    mem[14954] = 'd0;
    mem[14955] = 'd1020;
    mem[14956] = 'd0;
    mem[14957] = 'd0;
    mem[14958] = 'd0;
    mem[14959] = 'd1020;
    mem[14960] = 'd0;
    mem[14961] = 'd1020;
    mem[14962] = 'd0;
    mem[14963] = 'd0;
    mem[14964] = 'd0;
    mem[14965] = 'd1020;
    mem[14966] = 'd0;
    mem[14967] = 'd1020;
    mem[14968] = 'd0;
    mem[14969] = 'd0;
    mem[14970] = 'd0;
    mem[14971] = 'd1020;
    mem[14972] = 'd0;
    mem[14973] = 'd1020;
    mem[14974] = 'd0;
    mem[14975] = 'd0;
    mem[14976] = 'd0;
    mem[14977] = 'd0;
    mem[14978] = 'd1020;
    mem[14979] = 'd0;
    mem[14980] = 'd1020;
    mem[14981] = 'd0;
    mem[14982] = 'd0;
    mem[14983] = 'd0;
    mem[14984] = 'd1020;
    mem[14985] = 'd0;
    mem[14986] = 'd1020;
    mem[14987] = 'd0;
    mem[14988] = 'd0;
    mem[14989] = 'd0;
    mem[14990] = 'd1020;
    mem[14991] = 'd0;
    mem[14992] = 'd1020;
    mem[14993] = 'd0;
    mem[14994] = 'd0;
    mem[14995] = 'd0;
    mem[14996] = 'd1020;
    mem[14997] = 'd0;
    mem[14998] = 'd1020;
    mem[14999] = 'd0;
    mem[15000] = 'd0;
    mem[15001] = 'd0;
    mem[15002] = 'd1016;
    mem[15003] = 'd0;
    mem[15004] = 'd1020;
    mem[15005] = 'd0;
    mem[15006] = 'd0;
    mem[15007] = 'd0;
    mem[15008] = 'd1012;
    mem[15009] = 'd0;
    mem[15010] = 'd1020;
    mem[15011] = 'd0;
    mem[15012] = 'd0;
    mem[15013] = 'd0;
    mem[15014] = 'd896;
    mem[15015] = 'd0;
    mem[15016] = 'd940;
    mem[15017] = 'd0;
    mem[15018] = 'd0;
    mem[15019] = 'd0;
    mem[15020] = 'd220;
    mem[15021] = 'd0;
    mem[15022] = 'd540;
    mem[15023] = 'd0;
    mem[15024] = 'd0;
    mem[15025] = 'd0;
    mem[15026] = 'd20;
    mem[15027] = 'd0;
    mem[15028] = 'd476;
    mem[15029] = 'd0;
    mem[15030] = 'd0;
    mem[15031] = 'd0;
    mem[15032] = 'd36;
    mem[15033] = 'd0;
    mem[15034] = 'd528;
    mem[15035] = 'd0;
    mem[15036] = 'd0;
    mem[15037] = 'd0;
    mem[15038] = 'd52;
    mem[15039] = 'd0;
    mem[15040] = 'd572;
    mem[15041] = 'd0;
    mem[15042] = 'd0;
    mem[15043] = 'd0;
    mem[15044] = 'd64;
    mem[15045] = 'd0;
    mem[15046] = 'd600;
    mem[15047] = 'd0;
    mem[15048] = 'd0;
    mem[15049] = 'd0;
    mem[15050] = 'd72;
    mem[15051] = 'd0;
    mem[15052] = 'd624;
    mem[15053] = 'd0;
    mem[15054] = 'd0;
    mem[15055] = 'd0;
    mem[15056] = 'd80;
    mem[15057] = 'd0;
    mem[15058] = 'd640;
    mem[15059] = 'd0;
    mem[15060] = 'd0;
    mem[15061] = 'd0;
    mem[15062] = 'd84;
    mem[15063] = 'd0;
    mem[15064] = 'd656;
    mem[15065] = 'd0;
    mem[15066] = 'd0;
    mem[15067] = 'd0;
    mem[15068] = 'd88;
    mem[15069] = 'd0;
    mem[15070] = 'd664;
    mem[15071] = 'd0;
    mem[15072] = 'd0;
    mem[15073] = 'd0;
    mem[15074] = 'd88;
    mem[15075] = 'd0;
    mem[15076] = 'd668;
    mem[15077] = 'd0;
    mem[15078] = 'd0;
    mem[15079] = 'd0;
    mem[15080] = 'd92;
    mem[15081] = 'd0;
    mem[15082] = 'd672;
    mem[15083] = 'd0;
    mem[15084] = 'd0;
    mem[15085] = 'd0;
    mem[15086] = 'd88;
    mem[15087] = 'd0;
    mem[15088] = 'd672;
    mem[15089] = 'd0;
    mem[15090] = 'd0;
    mem[15091] = 'd0;
    mem[15092] = 'd88;
    mem[15093] = 'd0;
    mem[15094] = 'd672;
    mem[15095] = 'd0;
    mem[15096] = 'd0;
    mem[15097] = 'd0;
    mem[15098] = 'd88;
    mem[15099] = 'd0;
    mem[15100] = 'd672;
    mem[15101] = 'd0;
    mem[15102] = 'd0;
    mem[15103] = 'd0;
    mem[15104] = 'd88;
    mem[15105] = 'd0;
    mem[15106] = 'd668;
    mem[15107] = 'd0;
    mem[15108] = 'd0;
    mem[15109] = 'd0;
    mem[15110] = 'd88;
    mem[15111] = 'd0;
    mem[15112] = 'd664;
    mem[15113] = 'd0;
    mem[15114] = 'd0;
    mem[15115] = 'd0;
    mem[15116] = 'd84;
    mem[15117] = 'd0;
    mem[15118] = 'd656;
    mem[15119] = 'd0;
    mem[15120] = 'd0;
    mem[15121] = 'd0;
    mem[15122] = 'd80;
    mem[15123] = 'd0;
    mem[15124] = 'd644;
    mem[15125] = 'd0;
    mem[15126] = 'd0;
    mem[15127] = 'd0;
    mem[15128] = 'd72;
    mem[15129] = 'd0;
    mem[15130] = 'd628;
    mem[15131] = 'd0;
    mem[15132] = 'd0;
    mem[15133] = 'd0;
    mem[15134] = 'd64;
    mem[15135] = 'd0;
    mem[15136] = 'd604;
    mem[15137] = 'd0;
    mem[15138] = 'd0;
    mem[15139] = 'd0;
    mem[15140] = 'd56;
    mem[15141] = 'd0;
    mem[15142] = 'd572;
    mem[15143] = 'd0;
    mem[15144] = 'd0;
    mem[15145] = 'd0;
    mem[15146] = 'd36;
    mem[15147] = 'd0;
    mem[15148] = 'd532;
    mem[15149] = 'd0;
    mem[15150] = 'd0;
    mem[15151] = 'd0;
    mem[15152] = 'd24;
    mem[15153] = 'd0;
    mem[15154] = 'd480;
    mem[15155] = 'd0;
    mem[15156] = 'd0;
    mem[15157] = 'd0;
    mem[15158] = 'd196;
    mem[15159] = 'd0;
    mem[15160] = 'd520;
    mem[15161] = 'd0;
    mem[15162] = 'd0;
    mem[15163] = 'd0;
    mem[15164] = 'd892;
    mem[15165] = 'd0;
    mem[15166] = 'd940;
    mem[15167] = 'd0;
    mem[15168] = 'd0;
    mem[15169] = 'd0;
    mem[15170] = 'd1012;
    mem[15171] = 'd0;
    mem[15172] = 'd1016;
    mem[15173] = 'd0;
    mem[15174] = 'd0;
    mem[15175] = 'd0;
    mem[15176] = 'd1016;
    mem[15177] = 'd0;
    mem[15178] = 'd1020;
    mem[15179] = 'd0;
    mem[15180] = 'd0;
    mem[15181] = 'd0;
    mem[15182] = 'd1020;
    mem[15183] = 'd0;
    mem[15184] = 'd1020;
    mem[15185] = 'd0;
    mem[15186] = 'd0;
    mem[15187] = 'd0;
    mem[15188] = 'd1020;
    mem[15189] = 'd0;
    mem[15190] = 'd1020;
    mem[15191] = 'd0;
    mem[15192] = 'd0;
    mem[15193] = 'd0;
    mem[15194] = 'd1020;
    mem[15195] = 'd0;
    mem[15196] = 'd1020;
    mem[15197] = 'd0;
    mem[15198] = 'd0;
    mem[15199] = 'd0;
    mem[15200] = 'd1020;
    mem[15201] = 'd0;
    mem[15202] = 'd1020;
    mem[15203] = 'd0;
    mem[15204] = 'd0;
    mem[15205] = 'd0;
    mem[15206] = 'd1020;
    mem[15207] = 'd0;
    mem[15208] = 'd1020;
    mem[15209] = 'd0;
    mem[15210] = 'd0;
    mem[15211] = 'd1020;
    mem[15212] = 'd0;
    mem[15213] = 'd1020;
    mem[15214] = 'd0;
    mem[15215] = 'd0;
    mem[15216] = 'd0;
    mem[15217] = 'd1020;
    mem[15218] = 'd0;
    mem[15219] = 'd1020;
    mem[15220] = 'd0;
    mem[15221] = 'd0;
    mem[15222] = 'd0;
    mem[15223] = 'd1020;
    mem[15224] = 'd0;
    mem[15225] = 'd1020;
    mem[15226] = 'd0;
    mem[15227] = 'd0;
    mem[15228] = 'd0;
    mem[15229] = 'd1020;
    mem[15230] = 'd0;
    mem[15231] = 'd1020;
    mem[15232] = 'd0;
    mem[15233] = 'd0;
    mem[15234] = 'd0;
    mem[15235] = 'd1020;
    mem[15236] = 'd0;
    mem[15237] = 'd1020;
    mem[15238] = 'd0;
    mem[15239] = 'd0;
    mem[15240] = 'd0;
    mem[15241] = 'd1020;
    mem[15242] = 'd0;
    mem[15243] = 'd1020;
    mem[15244] = 'd0;
    mem[15245] = 'd0;
    mem[15246] = 'd0;
    mem[15247] = 'd940;
    mem[15248] = 'd0;
    mem[15249] = 'd988;
    mem[15250] = 'd0;
    mem[15251] = 'd0;
    mem[15252] = 'd0;
    mem[15253] = 'd540;
    mem[15254] = 'd0;
    mem[15255] = 'd840;
    mem[15256] = 'd0;
    mem[15257] = 'd0;
    mem[15258] = 'd0;
    mem[15259] = 'd476;
    mem[15260] = 'd0;
    mem[15261] = 'd844;
    mem[15262] = 'd0;
    mem[15263] = 'd0;
    mem[15264] = 'd0;
    mem[15265] = 'd528;
    mem[15266] = 'd0;
    mem[15267] = 'd876;
    mem[15268] = 'd0;
    mem[15269] = 'd0;
    mem[15270] = 'd0;
    mem[15271] = 'd572;
    mem[15272] = 'd0;
    mem[15273] = 'd900;
    mem[15274] = 'd0;
    mem[15275] = 'd0;
    mem[15276] = 'd0;
    mem[15277] = 'd600;
    mem[15278] = 'd0;
    mem[15279] = 'd924;
    mem[15280] = 'd0;
    mem[15281] = 'd0;
    mem[15282] = 'd0;
    mem[15283] = 'd624;
    mem[15284] = 'd0;
    mem[15285] = 'd948;
    mem[15286] = 'd0;
    mem[15287] = 'd0;
    mem[15288] = 'd0;
    mem[15289] = 'd640;
    mem[15290] = 'd0;
    mem[15291] = 'd964;
    mem[15292] = 'd0;
    mem[15293] = 'd0;
    mem[15294] = 'd0;
    mem[15295] = 'd656;
    mem[15296] = 'd0;
    mem[15297] = 'd980;
    mem[15298] = 'd0;
    mem[15299] = 'd0;
    mem[15300] = 'd0;
    mem[15301] = 'd664;
    mem[15302] = 'd0;
    mem[15303] = 'd988;
    mem[15304] = 'd0;
    mem[15305] = 'd0;
    mem[15306] = 'd0;
    mem[15307] = 'd668;
    mem[15308] = 'd0;
    mem[15309] = 'd996;
    mem[15310] = 'd0;
    mem[15311] = 'd0;
    mem[15312] = 'd0;
    mem[15313] = 'd672;
    mem[15314] = 'd0;
    mem[15315] = 'd996;
    mem[15316] = 'd0;
    mem[15317] = 'd0;
    mem[15318] = 'd0;
    mem[15319] = 'd672;
    mem[15320] = 'd0;
    mem[15321] = 'd1000;
    mem[15322] = 'd0;
    mem[15323] = 'd0;
    mem[15324] = 'd0;
    mem[15325] = 'd672;
    mem[15326] = 'd0;
    mem[15327] = 'd1000;
    mem[15328] = 'd0;
    mem[15329] = 'd0;
    mem[15330] = 'd0;
    mem[15331] = 'd672;
    mem[15332] = 'd0;
    mem[15333] = 'd996;
    mem[15334] = 'd0;
    mem[15335] = 'd0;
    mem[15336] = 'd0;
    mem[15337] = 'd668;
    mem[15338] = 'd0;
    mem[15339] = 'd996;
    mem[15340] = 'd0;
    mem[15341] = 'd0;
    mem[15342] = 'd0;
    mem[15343] = 'd664;
    mem[15344] = 'd0;
    mem[15345] = 'd988;
    mem[15346] = 'd0;
    mem[15347] = 'd0;
    mem[15348] = 'd0;
    mem[15349] = 'd656;
    mem[15350] = 'd0;
    mem[15351] = 'd980;
    mem[15352] = 'd0;
    mem[15353] = 'd0;
    mem[15354] = 'd0;
    mem[15355] = 'd644;
    mem[15356] = 'd0;
    mem[15357] = 'd964;
    mem[15358] = 'd0;
    mem[15359] = 'd0;
    mem[15360] = 'd0;
    mem[15361] = 'd628;
    mem[15362] = 'd0;
    mem[15363] = 'd948;
    mem[15364] = 'd0;
    mem[15365] = 'd0;
    mem[15366] = 'd0;
    mem[15367] = 'd604;
    mem[15368] = 'd0;
    mem[15369] = 'd928;
    mem[15370] = 'd0;
    mem[15371] = 'd0;
    mem[15372] = 'd0;
    mem[15373] = 'd572;
    mem[15374] = 'd0;
    mem[15375] = 'd904;
    mem[15376] = 'd0;
    mem[15377] = 'd0;
    mem[15378] = 'd0;
    mem[15379] = 'd532;
    mem[15380] = 'd0;
    mem[15381] = 'd880;
    mem[15382] = 'd0;
    mem[15383] = 'd0;
    mem[15384] = 'd0;
    mem[15385] = 'd480;
    mem[15386] = 'd0;
    mem[15387] = 'd848;
    mem[15388] = 'd0;
    mem[15389] = 'd0;
    mem[15390] = 'd0;
    mem[15391] = 'd520;
    mem[15392] = 'd0;
    mem[15393] = 'd832;
    mem[15394] = 'd0;
    mem[15395] = 'd0;
    mem[15396] = 'd0;
    mem[15397] = 'd940;
    mem[15398] = 'd0;
    mem[15399] = 'd988;
    mem[15400] = 'd0;
    mem[15401] = 'd0;
    mem[15402] = 'd0;
    mem[15403] = 'd1016;
    mem[15404] = 'd0;
    mem[15405] = 'd1020;
    mem[15406] = 'd0;
    mem[15407] = 'd0;
    mem[15408] = 'd0;
    mem[15409] = 'd1020;
    mem[15410] = 'd0;
    mem[15411] = 'd1020;
    mem[15412] = 'd0;
    mem[15413] = 'd0;
    mem[15414] = 'd0;
    mem[15415] = 'd1020;
    mem[15416] = 'd0;
    mem[15417] = 'd1020;
    mem[15418] = 'd0;
    mem[15419] = 'd0;
    mem[15420] = 'd0;
    mem[15421] = 'd1020;
    mem[15422] = 'd0;
    mem[15423] = 'd1020;
    mem[15424] = 'd0;
    mem[15425] = 'd0;
    mem[15426] = 'd0;
    mem[15427] = 'd1020;
    mem[15428] = 'd0;
    mem[15429] = 'd1020;
    mem[15430] = 'd0;
    mem[15431] = 'd0;
    mem[15432] = 'd0;
    mem[15433] = 'd1020;
    mem[15434] = 'd0;
    mem[15435] = 'd1020;
    mem[15436] = 'd0;
    mem[15437] = 'd0;
    mem[15438] = 'd0;
    mem[15439] = 'd1020;
    mem[15440] = 'd0;
    mem[15441] = 'd1020;
    mem[15442] = 'd0;
    mem[15443] = 'd0;
    mem[15444] = 'd0;
    mem[15445] = 'd0;
    mem[15446] = 'd1020;
    mem[15447] = 'd0;
    mem[15448] = 'd1020;
    mem[15449] = 'd0;
    mem[15450] = 'd0;
    mem[15451] = 'd0;
    mem[15452] = 'd1020;
    mem[15453] = 'd0;
    mem[15454] = 'd1020;
    mem[15455] = 'd0;
    mem[15456] = 'd0;
    mem[15457] = 'd0;
    mem[15458] = 'd1020;
    mem[15459] = 'd0;
    mem[15460] = 'd1020;
    mem[15461] = 'd0;
    mem[15462] = 'd0;
    mem[15463] = 'd0;
    mem[15464] = 'd1020;
    mem[15465] = 'd0;
    mem[15466] = 'd1020;
    mem[15467] = 'd0;
    mem[15468] = 'd0;
    mem[15469] = 'd0;
    mem[15470] = 'd1020;
    mem[15471] = 'd0;
    mem[15472] = 'd1020;
    mem[15473] = 'd0;
    mem[15474] = 'd0;
    mem[15475] = 'd0;
    mem[15476] = 'd1016;
    mem[15477] = 'd0;
    mem[15478] = 'd1020;
    mem[15479] = 'd0;
    mem[15480] = 'd0;
    mem[15481] = 'd0;
    mem[15482] = 'd1012;
    mem[15483] = 'd0;
    mem[15484] = 'd1020;
    mem[15485] = 'd0;
    mem[15486] = 'd0;
    mem[15487] = 'd0;
    mem[15488] = 'd944;
    mem[15489] = 'd0;
    mem[15490] = 'd976;
    mem[15491] = 'd0;
    mem[15492] = 'd0;
    mem[15493] = 'd0;
    mem[15494] = 'd416;
    mem[15495] = 'd0;
    mem[15496] = 'd664;
    mem[15497] = 'd0;
    mem[15498] = 'd0;
    mem[15499] = 'd0;
    mem[15500] = 'd24;
    mem[15501] = 'd0;
    mem[15502] = 'd456;
    mem[15503] = 'd0;
    mem[15504] = 'd0;
    mem[15505] = 'd0;
    mem[15506] = 'd28;
    mem[15507] = 'd0;
    mem[15508] = 'd504;
    mem[15509] = 'd0;
    mem[15510] = 'd0;
    mem[15511] = 'd0;
    mem[15512] = 'd40;
    mem[15513] = 'd0;
    mem[15514] = 'd544;
    mem[15515] = 'd0;
    mem[15516] = 'd0;
    mem[15517] = 'd0;
    mem[15518] = 'd52;
    mem[15519] = 'd0;
    mem[15520] = 'd576;
    mem[15521] = 'd0;
    mem[15522] = 'd0;
    mem[15523] = 'd0;
    mem[15524] = 'd60;
    mem[15525] = 'd0;
    mem[15526] = 'd596;
    mem[15527] = 'd0;
    mem[15528] = 'd0;
    mem[15529] = 'd0;
    mem[15530] = 'd68;
    mem[15531] = 'd0;
    mem[15532] = 'd616;
    mem[15533] = 'd0;
    mem[15534] = 'd0;
    mem[15535] = 'd0;
    mem[15536] = 'd72;
    mem[15537] = 'd0;
    mem[15538] = 'd628;
    mem[15539] = 'd0;
    mem[15540] = 'd0;
    mem[15541] = 'd0;
    mem[15542] = 'd76;
    mem[15543] = 'd0;
    mem[15544] = 'd636;
    mem[15545] = 'd0;
    mem[15546] = 'd0;
    mem[15547] = 'd0;
    mem[15548] = 'd80;
    mem[15549] = 'd0;
    mem[15550] = 'd644;
    mem[15551] = 'd0;
    mem[15552] = 'd0;
    mem[15553] = 'd0;
    mem[15554] = 'd80;
    mem[15555] = 'd0;
    mem[15556] = 'd644;
    mem[15557] = 'd0;
    mem[15558] = 'd0;
    mem[15559] = 'd0;
    mem[15560] = 'd80;
    mem[15561] = 'd0;
    mem[15562] = 'd644;
    mem[15563] = 'd0;
    mem[15564] = 'd0;
    mem[15565] = 'd0;
    mem[15566] = 'd80;
    mem[15567] = 'd0;
    mem[15568] = 'd640;
    mem[15569] = 'd0;
    mem[15570] = 'd0;
    mem[15571] = 'd0;
    mem[15572] = 'd76;
    mem[15573] = 'd0;
    mem[15574] = 'd636;
    mem[15575] = 'd0;
    mem[15576] = 'd0;
    mem[15577] = 'd0;
    mem[15578] = 'd72;
    mem[15579] = 'd0;
    mem[15580] = 'd628;
    mem[15581] = 'd0;
    mem[15582] = 'd0;
    mem[15583] = 'd0;
    mem[15584] = 'd68;
    mem[15585] = 'd0;
    mem[15586] = 'd620;
    mem[15587] = 'd0;
    mem[15588] = 'd0;
    mem[15589] = 'd0;
    mem[15590] = 'd60;
    mem[15591] = 'd0;
    mem[15592] = 'd600;
    mem[15593] = 'd0;
    mem[15594] = 'd0;
    mem[15595] = 'd0;
    mem[15596] = 'd52;
    mem[15597] = 'd0;
    mem[15598] = 'd580;
    mem[15599] = 'd0;
    mem[15600] = 'd0;
    mem[15601] = 'd0;
    mem[15602] = 'd44;
    mem[15603] = 'd0;
    mem[15604] = 'd548;
    mem[15605] = 'd0;
    mem[15606] = 'd0;
    mem[15607] = 'd0;
    mem[15608] = 'd32;
    mem[15609] = 'd0;
    mem[15610] = 'd508;
    mem[15611] = 'd0;
    mem[15612] = 'd0;
    mem[15613] = 'd0;
    mem[15614] = 'd24;
    mem[15615] = 'd0;
    mem[15616] = 'd456;
    mem[15617] = 'd0;
    mem[15618] = 'd0;
    mem[15619] = 'd0;
    mem[15620] = 'd388;
    mem[15621] = 'd0;
    mem[15622] = 'd648;
    mem[15623] = 'd0;
    mem[15624] = 'd0;
    mem[15625] = 'd0;
    mem[15626] = 'd932;
    mem[15627] = 'd0;
    mem[15628] = 'd968;
    mem[15629] = 'd0;
    mem[15630] = 'd0;
    mem[15631] = 'd0;
    mem[15632] = 'd1012;
    mem[15633] = 'd0;
    mem[15634] = 'd1016;
    mem[15635] = 'd0;
    mem[15636] = 'd0;
    mem[15637] = 'd0;
    mem[15638] = 'd1016;
    mem[15639] = 'd0;
    mem[15640] = 'd1020;
    mem[15641] = 'd0;
    mem[15642] = 'd0;
    mem[15643] = 'd0;
    mem[15644] = 'd1020;
    mem[15645] = 'd0;
    mem[15646] = 'd1020;
    mem[15647] = 'd0;
    mem[15648] = 'd0;
    mem[15649] = 'd0;
    mem[15650] = 'd1020;
    mem[15651] = 'd0;
    mem[15652] = 'd1020;
    mem[15653] = 'd0;
    mem[15654] = 'd0;
    mem[15655] = 'd0;
    mem[15656] = 'd1020;
    mem[15657] = 'd0;
    mem[15658] = 'd1020;
    mem[15659] = 'd0;
    mem[15660] = 'd0;
    mem[15661] = 'd0;
    mem[15662] = 'd1020;
    mem[15663] = 'd0;
    mem[15664] = 'd1020;
    mem[15665] = 'd0;
    mem[15666] = 'd0;
    mem[15667] = 'd0;
    mem[15668] = 'd1020;
    mem[15669] = 'd0;
    mem[15670] = 'd1020;
    mem[15671] = 'd0;
    mem[15672] = 'd0;
    mem[15673] = 'd0;
    mem[15674] = 'd1020;
    mem[15675] = 'd0;
    mem[15676] = 'd1020;
    mem[15677] = 'd0;
    mem[15678] = 'd0;
    mem[15679] = 'd1020;
    mem[15680] = 'd0;
    mem[15681] = 'd1020;
    mem[15682] = 'd0;
    mem[15683] = 'd0;
    mem[15684] = 'd0;
    mem[15685] = 'd1020;
    mem[15686] = 'd0;
    mem[15687] = 'd1020;
    mem[15688] = 'd0;
    mem[15689] = 'd0;
    mem[15690] = 'd0;
    mem[15691] = 'd1020;
    mem[15692] = 'd0;
    mem[15693] = 'd1020;
    mem[15694] = 'd0;
    mem[15695] = 'd0;
    mem[15696] = 'd0;
    mem[15697] = 'd1020;
    mem[15698] = 'd0;
    mem[15699] = 'd1020;
    mem[15700] = 'd0;
    mem[15701] = 'd0;
    mem[15702] = 'd0;
    mem[15703] = 'd1020;
    mem[15704] = 'd0;
    mem[15705] = 'd1020;
    mem[15706] = 'd0;
    mem[15707] = 'd0;
    mem[15708] = 'd0;
    mem[15709] = 'd1020;
    mem[15710] = 'd0;
    mem[15711] = 'd1020;
    mem[15712] = 'd0;
    mem[15713] = 'd0;
    mem[15714] = 'd0;
    mem[15715] = 'd1020;
    mem[15716] = 'd0;
    mem[15717] = 'd1020;
    mem[15718] = 'd0;
    mem[15719] = 'd0;
    mem[15720] = 'd0;
    mem[15721] = 'd976;
    mem[15722] = 'd0;
    mem[15723] = 'd1000;
    mem[15724] = 'd0;
    mem[15725] = 'd0;
    mem[15726] = 'd0;
    mem[15727] = 'd664;
    mem[15728] = 'd0;
    mem[15729] = 'd888;
    mem[15730] = 'd0;
    mem[15731] = 'd0;
    mem[15732] = 'd0;
    mem[15733] = 'd456;
    mem[15734] = 'd0;
    mem[15735] = 'd824;
    mem[15736] = 'd0;
    mem[15737] = 'd0;
    mem[15738] = 'd0;
    mem[15739] = 'd504;
    mem[15740] = 'd0;
    mem[15741] = 'd864;
    mem[15742] = 'd0;
    mem[15743] = 'd0;
    mem[15744] = 'd0;
    mem[15745] = 'd544;
    mem[15746] = 'd0;
    mem[15747] = 'd888;
    mem[15748] = 'd0;
    mem[15749] = 'd0;
    mem[15750] = 'd0;
    mem[15751] = 'd576;
    mem[15752] = 'd0;
    mem[15753] = 'd908;
    mem[15754] = 'd0;
    mem[15755] = 'd0;
    mem[15756] = 'd0;
    mem[15757] = 'd596;
    mem[15758] = 'd0;
    mem[15759] = 'd924;
    mem[15760] = 'd0;
    mem[15761] = 'd0;
    mem[15762] = 'd0;
    mem[15763] = 'd616;
    mem[15764] = 'd0;
    mem[15765] = 'd944;
    mem[15766] = 'd0;
    mem[15767] = 'd0;
    mem[15768] = 'd0;
    mem[15769] = 'd628;
    mem[15770] = 'd0;
    mem[15771] = 'd952;
    mem[15772] = 'd0;
    mem[15773] = 'd0;
    mem[15774] = 'd0;
    mem[15775] = 'd636;
    mem[15776] = 'd0;
    mem[15777] = 'd964;
    mem[15778] = 'd0;
    mem[15779] = 'd0;
    mem[15780] = 'd0;
    mem[15781] = 'd644;
    mem[15782] = 'd0;
    mem[15783] = 'd964;
    mem[15784] = 'd0;
    mem[15785] = 'd0;
    mem[15786] = 'd0;
    mem[15787] = 'd644;
    mem[15788] = 'd0;
    mem[15789] = 'd968;
    mem[15790] = 'd0;
    mem[15791] = 'd0;
    mem[15792] = 'd0;
    mem[15793] = 'd644;
    mem[15794] = 'd0;
    mem[15795] = 'd968;
    mem[15796] = 'd0;
    mem[15797] = 'd0;
    mem[15798] = 'd0;
    mem[15799] = 'd640;
    mem[15800] = 'd0;
    mem[15801] = 'd968;
    mem[15802] = 'd0;
    mem[15803] = 'd0;
    mem[15804] = 'd0;
    mem[15805] = 'd636;
    mem[15806] = 'd0;
    mem[15807] = 'd964;
    mem[15808] = 'd0;
    mem[15809] = 'd0;
    mem[15810] = 'd0;
    mem[15811] = 'd628;
    mem[15812] = 'd0;
    mem[15813] = 'd956;
    mem[15814] = 'd0;
    mem[15815] = 'd0;
    mem[15816] = 'd0;
    mem[15817] = 'd620;
    mem[15818] = 'd0;
    mem[15819] = 'd944;
    mem[15820] = 'd0;
    mem[15821] = 'd0;
    mem[15822] = 'd0;
    mem[15823] = 'd600;
    mem[15824] = 'd0;
    mem[15825] = 'd928;
    mem[15826] = 'd0;
    mem[15827] = 'd0;
    mem[15828] = 'd0;
    mem[15829] = 'd580;
    mem[15830] = 'd0;
    mem[15831] = 'd912;
    mem[15832] = 'd0;
    mem[15833] = 'd0;
    mem[15834] = 'd0;
    mem[15835] = 'd548;
    mem[15836] = 'd0;
    mem[15837] = 'd892;
    mem[15838] = 'd0;
    mem[15839] = 'd0;
    mem[15840] = 'd0;
    mem[15841] = 'd508;
    mem[15842] = 'd0;
    mem[15843] = 'd868;
    mem[15844] = 'd0;
    mem[15845] = 'd0;
    mem[15846] = 'd0;
    mem[15847] = 'd456;
    mem[15848] = 'd0;
    mem[15849] = 'd828;
    mem[15850] = 'd0;
    mem[15851] = 'd0;
    mem[15852] = 'd0;
    mem[15853] = 'd648;
    mem[15854] = 'd0;
    mem[15855] = 'd884;
    mem[15856] = 'd0;
    mem[15857] = 'd0;
    mem[15858] = 'd0;
    mem[15859] = 'd968;
    mem[15860] = 'd0;
    mem[15861] = 'd1000;
    mem[15862] = 'd0;
    mem[15863] = 'd0;
    mem[15864] = 'd0;
    mem[15865] = 'd1016;
    mem[15866] = 'd0;
    mem[15867] = 'd1020;
    mem[15868] = 'd0;
    mem[15869] = 'd0;
    mem[15870] = 'd0;
    mem[15871] = 'd1020;
    mem[15872] = 'd0;
    mem[15873] = 'd1020;
    mem[15874] = 'd0;
    mem[15875] = 'd0;
    mem[15876] = 'd0;
    mem[15877] = 'd1020;
    mem[15878] = 'd0;
    mem[15879] = 'd1020;
    mem[15880] = 'd0;
    mem[15881] = 'd0;
    mem[15882] = 'd0;
    mem[15883] = 'd1020;
    mem[15884] = 'd0;
    mem[15885] = 'd1020;
    mem[15886] = 'd0;
    mem[15887] = 'd0;
    mem[15888] = 'd0;
    mem[15889] = 'd1020;
    mem[15890] = 'd0;
    mem[15891] = 'd1020;
    mem[15892] = 'd0;
    mem[15893] = 'd0;
    mem[15894] = 'd0;
    mem[15895] = 'd1020;
    mem[15896] = 'd0;
    mem[15897] = 'd1020;
    mem[15898] = 'd0;
    mem[15899] = 'd0;
    mem[15900] = 'd0;
    mem[15901] = 'd1020;
    mem[15902] = 'd0;
    mem[15903] = 'd1020;
    mem[15904] = 'd0;
    mem[15905] = 'd0;
    mem[15906] = 'd0;
    mem[15907] = 'd1020;
    mem[15908] = 'd0;
    mem[15909] = 'd1020;
    mem[15910] = 'd0;
    mem[15911] = 'd0;
    mem[15912] = 'd0;
    mem[15913] = 'd0;
    mem[15914] = 'd1020;
    mem[15915] = 'd0;
    mem[15916] = 'd1020;
    mem[15917] = 'd0;
    mem[15918] = 'd0;
    mem[15919] = 'd0;
    mem[15920] = 'd1020;
    mem[15921] = 'd0;
    mem[15922] = 'd1020;
    mem[15923] = 'd0;
    mem[15924] = 'd0;
    mem[15925] = 'd0;
    mem[15926] = 'd1020;
    mem[15927] = 'd0;
    mem[15928] = 'd1020;
    mem[15929] = 'd0;
    mem[15930] = 'd0;
    mem[15931] = 'd0;
    mem[15932] = 'd1020;
    mem[15933] = 'd0;
    mem[15934] = 'd1020;
    mem[15935] = 'd0;
    mem[15936] = 'd0;
    mem[15937] = 'd0;
    mem[15938] = 'd1020;
    mem[15939] = 'd0;
    mem[15940] = 'd1020;
    mem[15941] = 'd0;
    mem[15942] = 'd0;
    mem[15943] = 'd0;
    mem[15944] = 'd1020;
    mem[15945] = 'd0;
    mem[15946] = 'd1020;
    mem[15947] = 'd0;
    mem[15948] = 'd0;
    mem[15949] = 'd0;
    mem[15950] = 'd1016;
    mem[15951] = 'd0;
    mem[15952] = 'd1020;
    mem[15953] = 'd0;
    mem[15954] = 'd0;
    mem[15955] = 'd0;
    mem[15956] = 'd1012;
    mem[15957] = 'd0;
    mem[15958] = 'd1020;
    mem[15959] = 'd0;
    mem[15960] = 'd0;
    mem[15961] = 'd0;
    mem[15962] = 'd1004;
    mem[15963] = 'd0;
    mem[15964] = 'd1012;
    mem[15965] = 'd0;
    mem[15966] = 'd0;
    mem[15967] = 'd0;
    mem[15968] = 'd708;
    mem[15969] = 'd0;
    mem[15970] = 'd832;
    mem[15971] = 'd0;
    mem[15972] = 'd0;
    mem[15973] = 'd0;
    mem[15974] = 'd180;
    mem[15975] = 'd0;
    mem[15976] = 'd520;
    mem[15977] = 'd0;
    mem[15978] = 'd0;
    mem[15979] = 'd0;
    mem[15980] = 'd16;
    mem[15981] = 'd0;
    mem[15982] = 'd460;
    mem[15983] = 'd0;
    mem[15984] = 'd0;
    mem[15985] = 'd0;
    mem[15986] = 'd28;
    mem[15987] = 'd0;
    mem[15988] = 'd508;
    mem[15989] = 'd0;
    mem[15990] = 'd0;
    mem[15991] = 'd0;
    mem[15992] = 'd40;
    mem[15993] = 'd0;
    mem[15994] = 'd536;
    mem[15995] = 'd0;
    mem[15996] = 'd0;
    mem[15997] = 'd0;
    mem[15998] = 'd48;
    mem[15999] = 'd0;
    mem[16000] = 'd560;
    mem[16001] = 'd0;
    mem[16002] = 'd0;
    mem[16003] = 'd0;
    mem[16004] = 'd52;
    mem[16005] = 'd0;
    mem[16006] = 'd580;
    mem[16007] = 'd0;
    mem[16008] = 'd0;
    mem[16009] = 'd0;
    mem[16010] = 'd56;
    mem[16011] = 'd0;
    mem[16012] = 'd588;
    mem[16013] = 'd0;
    mem[16014] = 'd0;
    mem[16015] = 'd0;
    mem[16016] = 'd60;
    mem[16017] = 'd0;
    mem[16018] = 'd596;
    mem[16019] = 'd0;
    mem[16020] = 'd0;
    mem[16021] = 'd0;
    mem[16022] = 'd60;
    mem[16023] = 'd0;
    mem[16024] = 'd600;
    mem[16025] = 'd0;
    mem[16026] = 'd0;
    mem[16027] = 'd0;
    mem[16028] = 'd60;
    mem[16029] = 'd0;
    mem[16030] = 'd600;
    mem[16031] = 'd0;
    mem[16032] = 'd0;
    mem[16033] = 'd0;
    mem[16034] = 'd60;
    mem[16035] = 'd0;
    mem[16036] = 'd600;
    mem[16037] = 'd0;
    mem[16038] = 'd0;
    mem[16039] = 'd0;
    mem[16040] = 'd56;
    mem[16041] = 'd0;
    mem[16042] = 'd592;
    mem[16043] = 'd0;
    mem[16044] = 'd0;
    mem[16045] = 'd0;
    mem[16046] = 'd52;
    mem[16047] = 'd0;
    mem[16048] = 'd580;
    mem[16049] = 'd0;
    mem[16050] = 'd0;
    mem[16051] = 'd0;
    mem[16052] = 'd48;
    mem[16053] = 'd0;
    mem[16054] = 'd564;
    mem[16055] = 'd0;
    mem[16056] = 'd0;
    mem[16057] = 'd0;
    mem[16058] = 'd40;
    mem[16059] = 'd0;
    mem[16060] = 'd540;
    mem[16061] = 'd0;
    mem[16062] = 'd0;
    mem[16063] = 'd0;
    mem[16064] = 'd28;
    mem[16065] = 'd0;
    mem[16066] = 'd508;
    mem[16067] = 'd0;
    mem[16068] = 'd0;
    mem[16069] = 'd0;
    mem[16070] = 'd20;
    mem[16071] = 'd0;
    mem[16072] = 'd464;
    mem[16073] = 'd0;
    mem[16074] = 'd0;
    mem[16075] = 'd0;
    mem[16076] = 'd168;
    mem[16077] = 'd0;
    mem[16078] = 'd512;
    mem[16079] = 'd0;
    mem[16080] = 'd0;
    mem[16081] = 'd0;
    mem[16082] = 'd680;
    mem[16083] = 'd0;
    mem[16084] = 'd820;
    mem[16085] = 'd0;
    mem[16086] = 'd0;
    mem[16087] = 'd0;
    mem[16088] = 'd1000;
    mem[16089] = 'd0;
    mem[16090] = 'd1012;
    mem[16091] = 'd0;
    mem[16092] = 'd0;
    mem[16093] = 'd0;
    mem[16094] = 'd1012;
    mem[16095] = 'd0;
    mem[16096] = 'd1016;
    mem[16097] = 'd0;
    mem[16098] = 'd0;
    mem[16099] = 'd0;
    mem[16100] = 'd1016;
    mem[16101] = 'd0;
    mem[16102] = 'd1020;
    mem[16103] = 'd0;
    mem[16104] = 'd0;
    mem[16105] = 'd0;
    mem[16106] = 'd1020;
    mem[16107] = 'd0;
    mem[16108] = 'd1020;
    mem[16109] = 'd0;
    mem[16110] = 'd0;
    mem[16111] = 'd0;
    mem[16112] = 'd1020;
    mem[16113] = 'd0;
    mem[16114] = 'd1020;
    mem[16115] = 'd0;
    mem[16116] = 'd0;
    mem[16117] = 'd0;
    mem[16118] = 'd1020;
    mem[16119] = 'd0;
    mem[16120] = 'd1020;
    mem[16121] = 'd0;
    mem[16122] = 'd0;
    mem[16123] = 'd0;
    mem[16124] = 'd1020;
    mem[16125] = 'd0;
    mem[16126] = 'd1020;
    mem[16127] = 'd0;
    mem[16128] = 'd0;
    mem[16129] = 'd0;
    mem[16130] = 'd1020;
    mem[16131] = 'd0;
    mem[16132] = 'd1020;
    mem[16133] = 'd0;
    mem[16134] = 'd0;
    mem[16135] = 'd0;
    mem[16136] = 'd1020;
    mem[16137] = 'd0;
    mem[16138] = 'd1020;
    mem[16139] = 'd0;
    mem[16140] = 'd0;
    mem[16141] = 'd0;
    mem[16142] = 'd1020;
    mem[16143] = 'd0;
    mem[16144] = 'd1020;
    mem[16145] = 'd0;
    mem[16146] = 'd0;
    mem[16147] = 'd1020;
    mem[16148] = 'd0;
    mem[16149] = 'd1020;
    mem[16150] = 'd0;
    mem[16151] = 'd0;
    mem[16152] = 'd0;
    mem[16153] = 'd1020;
    mem[16154] = 'd0;
    mem[16155] = 'd1020;
    mem[16156] = 'd0;
    mem[16157] = 'd0;
    mem[16158] = 'd0;
    mem[16159] = 'd1020;
    mem[16160] = 'd0;
    mem[16161] = 'd1020;
    mem[16162] = 'd0;
    mem[16163] = 'd0;
    mem[16164] = 'd0;
    mem[16165] = 'd1020;
    mem[16166] = 'd0;
    mem[16167] = 'd1020;
    mem[16168] = 'd0;
    mem[16169] = 'd0;
    mem[16170] = 'd0;
    mem[16171] = 'd1020;
    mem[16172] = 'd0;
    mem[16173] = 'd1020;
    mem[16174] = 'd0;
    mem[16175] = 'd0;
    mem[16176] = 'd0;
    mem[16177] = 'd1020;
    mem[16178] = 'd0;
    mem[16179] = 'd1020;
    mem[16180] = 'd0;
    mem[16181] = 'd0;
    mem[16182] = 'd0;
    mem[16183] = 'd1020;
    mem[16184] = 'd0;
    mem[16185] = 'd1020;
    mem[16186] = 'd0;
    mem[16187] = 'd0;
    mem[16188] = 'd0;
    mem[16189] = 'd1020;
    mem[16190] = 'd0;
    mem[16191] = 'd1020;
    mem[16192] = 'd0;
    mem[16193] = 'd0;
    mem[16194] = 'd0;
    mem[16195] = 'd1012;
    mem[16196] = 'd0;
    mem[16197] = 'd1020;
    mem[16198] = 'd0;
    mem[16199] = 'd0;
    mem[16200] = 'd0;
    mem[16201] = 'd832;
    mem[16202] = 'd0;
    mem[16203] = 'd944;
    mem[16204] = 'd0;
    mem[16205] = 'd0;
    mem[16206] = 'd0;
    mem[16207] = 'd520;
    mem[16208] = 'd0;
    mem[16209] = 'd832;
    mem[16210] = 'd0;
    mem[16211] = 'd0;
    mem[16212] = 'd0;
    mem[16213] = 'd460;
    mem[16214] = 'd0;
    mem[16215] = 'd836;
    mem[16216] = 'd0;
    mem[16217] = 'd0;
    mem[16218] = 'd0;
    mem[16219] = 'd508;
    mem[16220] = 'd0;
    mem[16221] = 'd868;
    mem[16222] = 'd0;
    mem[16223] = 'd0;
    mem[16224] = 'd0;
    mem[16225] = 'd536;
    mem[16226] = 'd0;
    mem[16227] = 'd888;
    mem[16228] = 'd0;
    mem[16229] = 'd0;
    mem[16230] = 'd0;
    mem[16231] = 'd560;
    mem[16232] = 'd0;
    mem[16233] = 'd904;
    mem[16234] = 'd0;
    mem[16235] = 'd0;
    mem[16236] = 'd0;
    mem[16237] = 'd580;
    mem[16238] = 'd0;
    mem[16239] = 'd912;
    mem[16240] = 'd0;
    mem[16241] = 'd0;
    mem[16242] = 'd0;
    mem[16243] = 'd588;
    mem[16244] = 'd0;
    mem[16245] = 'd924;
    mem[16246] = 'd0;
    mem[16247] = 'd0;
    mem[16248] = 'd0;
    mem[16249] = 'd596;
    mem[16250] = 'd0;
    mem[16251] = 'd928;
    mem[16252] = 'd0;
    mem[16253] = 'd0;
    mem[16254] = 'd0;
    mem[16255] = 'd600;
    mem[16256] = 'd0;
    mem[16257] = 'd932;
    mem[16258] = 'd0;
    mem[16259] = 'd0;
    mem[16260] = 'd0;
    mem[16261] = 'd600;
    mem[16262] = 'd0;
    mem[16263] = 'd932;
    mem[16264] = 'd0;
    mem[16265] = 'd0;
    mem[16266] = 'd0;
    mem[16267] = 'd600;
    mem[16268] = 'd0;
    mem[16269] = 'd932;
    mem[16270] = 'd0;
    mem[16271] = 'd0;
    mem[16272] = 'd0;
    mem[16273] = 'd592;
    mem[16274] = 'd0;
    mem[16275] = 'd924;
    mem[16276] = 'd0;
    mem[16277] = 'd0;
    mem[16278] = 'd0;
    mem[16279] = 'd580;
    mem[16280] = 'd0;
    mem[16281] = 'd916;
    mem[16282] = 'd0;
    mem[16283] = 'd0;
    mem[16284] = 'd0;
    mem[16285] = 'd564;
    mem[16286] = 'd0;
    mem[16287] = 'd904;
    mem[16288] = 'd0;
    mem[16289] = 'd0;
    mem[16290] = 'd0;
    mem[16291] = 'd540;
    mem[16292] = 'd0;
    mem[16293] = 'd888;
    mem[16294] = 'd0;
    mem[16295] = 'd0;
    mem[16296] = 'd0;
    mem[16297] = 'd508;
    mem[16298] = 'd0;
    mem[16299] = 'd868;
    mem[16300] = 'd0;
    mem[16301] = 'd0;
    mem[16302] = 'd0;
    mem[16303] = 'd464;
    mem[16304] = 'd0;
    mem[16305] = 'd840;
    mem[16306] = 'd0;
    mem[16307] = 'd0;
    mem[16308] = 'd0;
    mem[16309] = 'd512;
    mem[16310] = 'd0;
    mem[16311] = 'd832;
    mem[16312] = 'd0;
    mem[16313] = 'd0;
    mem[16314] = 'd0;
    mem[16315] = 'd820;
    mem[16316] = 'd0;
    mem[16317] = 'd940;
    mem[16318] = 'd0;
    mem[16319] = 'd0;
    mem[16320] = 'd0;
    mem[16321] = 'd1012;
    mem[16322] = 'd0;
    mem[16323] = 'd1020;
    mem[16324] = 'd0;
    mem[16325] = 'd0;
    mem[16326] = 'd0;
    mem[16327] = 'd1016;
    mem[16328] = 'd0;
    mem[16329] = 'd1020;
    mem[16330] = 'd0;
    mem[16331] = 'd0;
    mem[16332] = 'd0;
    mem[16333] = 'd1020;
    mem[16334] = 'd0;
    mem[16335] = 'd1020;
    mem[16336] = 'd0;
    mem[16337] = 'd0;
    mem[16338] = 'd0;
    mem[16339] = 'd1020;
    mem[16340] = 'd0;
    mem[16341] = 'd1020;
    mem[16342] = 'd0;
    mem[16343] = 'd0;
    mem[16344] = 'd0;
    mem[16345] = 'd1020;
    mem[16346] = 'd0;
    mem[16347] = 'd1020;
    mem[16348] = 'd0;
    mem[16349] = 'd0;
    mem[16350] = 'd0;
    mem[16351] = 'd1020;
    mem[16352] = 'd0;
    mem[16353] = 'd1020;
    mem[16354] = 'd0;
    mem[16355] = 'd0;
    mem[16356] = 'd0;
    mem[16357] = 'd1020;
    mem[16358] = 'd0;
    mem[16359] = 'd1020;
    mem[16360] = 'd0;
    mem[16361] = 'd0;
    mem[16362] = 'd0;
    mem[16363] = 'd1020;
    mem[16364] = 'd0;
    mem[16365] = 'd1020;
    mem[16366] = 'd0;
    mem[16367] = 'd0;
    mem[16368] = 'd0;
    mem[16369] = 'd1020;
    mem[16370] = 'd0;
    mem[16371] = 'd1020;
    mem[16372] = 'd0;
    mem[16373] = 'd0;
    mem[16374] = 'd0;
    mem[16375] = 'd1020;
    mem[16376] = 'd0;
    mem[16377] = 'd1020;
    mem[16378] = 'd0;
    mem[16379] = 'd0;
    mem[16380] = 'd0;
    mem[16381] = 'd0;
    mem[16382] = 'd1020;
    mem[16383] = 'd0;
    mem[16384] = 'd1020;
    mem[16385] = 'd0;
    mem[16386] = 'd0;
    mem[16387] = 'd0;
    mem[16388] = 'd1020;
    mem[16389] = 'd0;
    mem[16390] = 'd1020;
    mem[16391] = 'd0;
    mem[16392] = 'd0;
    mem[16393] = 'd0;
    mem[16394] = 'd1020;
    mem[16395] = 'd0;
    mem[16396] = 'd1020;
    mem[16397] = 'd0;
    mem[16398] = 'd0;
    mem[16399] = 'd0;
    mem[16400] = 'd1020;
    mem[16401] = 'd0;
    mem[16402] = 'd1020;
    mem[16403] = 'd0;
    mem[16404] = 'd0;
    mem[16405] = 'd0;
    mem[16406] = 'd1020;
    mem[16407] = 'd0;
    mem[16408] = 'd1020;
    mem[16409] = 'd0;
    mem[16410] = 'd0;
    mem[16411] = 'd0;
    mem[16412] = 'd1020;
    mem[16413] = 'd0;
    mem[16414] = 'd1020;
    mem[16415] = 'd0;
    mem[16416] = 'd0;
    mem[16417] = 'd0;
    mem[16418] = 'd1020;
    mem[16419] = 'd0;
    mem[16420] = 'd1020;
    mem[16421] = 'd0;
    mem[16422] = 'd0;
    mem[16423] = 'd0;
    mem[16424] = 'd1020;
    mem[16425] = 'd0;
    mem[16426] = 'd1020;
    mem[16427] = 'd0;
    mem[16428] = 'd0;
    mem[16429] = 'd0;
    mem[16430] = 'd1016;
    mem[16431] = 'd0;
    mem[16432] = 'd1020;
    mem[16433] = 'd0;
    mem[16434] = 'd0;
    mem[16435] = 'd0;
    mem[16436] = 'd1008;
    mem[16437] = 'd0;
    mem[16438] = 'd1016;
    mem[16439] = 'd0;
    mem[16440] = 'd0;
    mem[16441] = 'd0;
    mem[16442] = 'd968;
    mem[16443] = 'd0;
    mem[16444] = 'd992;
    mem[16445] = 'd0;
    mem[16446] = 'd0;
    mem[16447] = 'd0;
    mem[16448] = 'd724;
    mem[16449] = 'd0;
    mem[16450] = 'd840;
    mem[16451] = 'd0;
    mem[16452] = 'd0;
    mem[16453] = 'd0;
    mem[16454] = 'd336;
    mem[16455] = 'd0;
    mem[16456] = 'd604;
    mem[16457] = 'd0;
    mem[16458] = 'd0;
    mem[16459] = 'd0;
    mem[16460] = 'd68;
    mem[16461] = 'd0;
    mem[16462] = 'd464;
    mem[16463] = 'd0;
    mem[16464] = 'd0;
    mem[16465] = 'd0;
    mem[16466] = 'd16;
    mem[16467] = 'd0;
    mem[16468] = 'd468;
    mem[16469] = 'd0;
    mem[16470] = 'd0;
    mem[16471] = 'd0;
    mem[16472] = 'd24;
    mem[16473] = 'd0;
    mem[16474] = 'd496;
    mem[16475] = 'd0;
    mem[16476] = 'd0;
    mem[16477] = 'd0;
    mem[16478] = 'd28;
    mem[16479] = 'd0;
    mem[16480] = 'd512;
    mem[16481] = 'd0;
    mem[16482] = 'd0;
    mem[16483] = 'd0;
    mem[16484] = 'd32;
    mem[16485] = 'd0;
    mem[16486] = 'd524;
    mem[16487] = 'd0;
    mem[16488] = 'd0;
    mem[16489] = 'd0;
    mem[16490] = 'd32;
    mem[16491] = 'd0;
    mem[16492] = 'd528;
    mem[16493] = 'd0;
    mem[16494] = 'd0;
    mem[16495] = 'd0;
    mem[16496] = 'd32;
    mem[16497] = 'd0;
    mem[16498] = 'd528;
    mem[16499] = 'd0;
    mem[16500] = 'd0;
    mem[16501] = 'd0;
    mem[16502] = 'd32;
    mem[16503] = 'd0;
    mem[16504] = 'd524;
    mem[16505] = 'd0;
    mem[16506] = 'd0;
    mem[16507] = 'd0;
    mem[16508] = 'd32;
    mem[16509] = 'd0;
    mem[16510] = 'd512;
    mem[16511] = 'd0;
    mem[16512] = 'd0;
    mem[16513] = 'd0;
    mem[16514] = 'd24;
    mem[16515] = 'd0;
    mem[16516] = 'd496;
    mem[16517] = 'd0;
    mem[16518] = 'd0;
    mem[16519] = 'd0;
    mem[16520] = 'd20;
    mem[16521] = 'd0;
    mem[16522] = 'd472;
    mem[16523] = 'd0;
    mem[16524] = 'd0;
    mem[16525] = 'd0;
    mem[16526] = 'd32;
    mem[16527] = 'd0;
    mem[16528] = 'd436;
    mem[16529] = 'd0;
    mem[16530] = 'd0;
    mem[16531] = 'd0;
    mem[16532] = 'd328;
    mem[16533] = 'd0;
    mem[16534] = 'd608;
    mem[16535] = 'd0;
    mem[16536] = 'd0;
    mem[16537] = 'd0;
    mem[16538] = 'd720;
    mem[16539] = 'd0;
    mem[16540] = 'd836;
    mem[16541] = 'd0;
    mem[16542] = 'd0;
    mem[16543] = 'd0;
    mem[16544] = 'd972;
    mem[16545] = 'd0;
    mem[16546] = 'd996;
    mem[16547] = 'd0;
    mem[16548] = 'd0;
    mem[16549] = 'd0;
    mem[16550] = 'd1008;
    mem[16551] = 'd0;
    mem[16552] = 'd1016;
    mem[16553] = 'd0;
    mem[16554] = 'd0;
    mem[16555] = 'd0;
    mem[16556] = 'd1012;
    mem[16557] = 'd0;
    mem[16558] = 'd1020;
    mem[16559] = 'd0;
    mem[16560] = 'd0;
    mem[16561] = 'd0;
    mem[16562] = 'd1016;
    mem[16563] = 'd0;
    mem[16564] = 'd1020;
    mem[16565] = 'd0;
    mem[16566] = 'd0;
    mem[16567] = 'd0;
    mem[16568] = 'd1020;
    mem[16569] = 'd0;
    mem[16570] = 'd1020;
    mem[16571] = 'd0;
    mem[16572] = 'd0;
    mem[16573] = 'd0;
    mem[16574] = 'd1020;
    mem[16575] = 'd0;
    mem[16576] = 'd1020;
    mem[16577] = 'd0;
    mem[16578] = 'd0;
    mem[16579] = 'd0;
    mem[16580] = 'd1020;
    mem[16581] = 'd0;
    mem[16582] = 'd1020;
    mem[16583] = 'd0;
    mem[16584] = 'd0;
    mem[16585] = 'd0;
    mem[16586] = 'd1020;
    mem[16587] = 'd0;
    mem[16588] = 'd1020;
    mem[16589] = 'd0;
    mem[16590] = 'd0;
    mem[16591] = 'd0;
    mem[16592] = 'd1020;
    mem[16593] = 'd0;
    mem[16594] = 'd1020;
    mem[16595] = 'd0;
    mem[16596] = 'd0;
    mem[16597] = 'd0;
    mem[16598] = 'd1020;
    mem[16599] = 'd0;
    mem[16600] = 'd1020;
    mem[16601] = 'd0;
    mem[16602] = 'd0;
    mem[16603] = 'd0;
    mem[16604] = 'd1020;
    mem[16605] = 'd0;
    mem[16606] = 'd1020;
    mem[16607] = 'd0;
    mem[16608] = 'd0;
    mem[16609] = 'd0;
    mem[16610] = 'd1020;
    mem[16611] = 'd0;
    mem[16612] = 'd1020;
    mem[16613] = 'd0;
    mem[16614] = 'd0;
    mem[16615] = 'd1020;
    mem[16616] = 'd0;
    mem[16617] = 'd1020;
    mem[16618] = 'd0;
    mem[16619] = 'd0;
    mem[16620] = 'd0;
    mem[16621] = 'd1020;
    mem[16622] = 'd0;
    mem[16623] = 'd1020;
    mem[16624] = 'd0;
    mem[16625] = 'd0;
    mem[16626] = 'd0;
    mem[16627] = 'd1020;
    mem[16628] = 'd0;
    mem[16629] = 'd1020;
    mem[16630] = 'd0;
    mem[16631] = 'd0;
    mem[16632] = 'd0;
    mem[16633] = 'd1020;
    mem[16634] = 'd0;
    mem[16635] = 'd1020;
    mem[16636] = 'd0;
    mem[16637] = 'd0;
    mem[16638] = 'd0;
    mem[16639] = 'd1020;
    mem[16640] = 'd0;
    mem[16641] = 'd1020;
    mem[16642] = 'd0;
    mem[16643] = 'd0;
    mem[16644] = 'd0;
    mem[16645] = 'd1020;
    mem[16646] = 'd0;
    mem[16647] = 'd1020;
    mem[16648] = 'd0;
    mem[16649] = 'd0;
    mem[16650] = 'd0;
    mem[16651] = 'd1020;
    mem[16652] = 'd0;
    mem[16653] = 'd1020;
    mem[16654] = 'd0;
    mem[16655] = 'd0;
    mem[16656] = 'd0;
    mem[16657] = 'd1020;
    mem[16658] = 'd0;
    mem[16659] = 'd1020;
    mem[16660] = 'd0;
    mem[16661] = 'd0;
    mem[16662] = 'd0;
    mem[16663] = 'd1020;
    mem[16664] = 'd0;
    mem[16665] = 'd1020;
    mem[16666] = 'd0;
    mem[16667] = 'd0;
    mem[16668] = 'd0;
    mem[16669] = 'd1016;
    mem[16670] = 'd0;
    mem[16671] = 'd1020;
    mem[16672] = 'd0;
    mem[16673] = 'd0;
    mem[16674] = 'd0;
    mem[16675] = 'd992;
    mem[16676] = 'd0;
    mem[16677] = 'd1008;
    mem[16678] = 'd0;
    mem[16679] = 'd0;
    mem[16680] = 'd0;
    mem[16681] = 'd840;
    mem[16682] = 'd0;
    mem[16683] = 'd952;
    mem[16684] = 'd0;
    mem[16685] = 'd0;
    mem[16686] = 'd0;
    mem[16687] = 'd604;
    mem[16688] = 'd0;
    mem[16689] = 'd856;
    mem[16690] = 'd0;
    mem[16691] = 'd0;
    mem[16692] = 'd0;
    mem[16693] = 'd464;
    mem[16694] = 'd0;
    mem[16695] = 'd816;
    mem[16696] = 'd0;
    mem[16697] = 'd0;
    mem[16698] = 'd0;
    mem[16699] = 'd468;
    mem[16700] = 'd0;
    mem[16701] = 'd840;
    mem[16702] = 'd0;
    mem[16703] = 'd0;
    mem[16704] = 'd0;
    mem[16705] = 'd496;
    mem[16706] = 'd0;
    mem[16707] = 'd860;
    mem[16708] = 'd0;
    mem[16709] = 'd0;
    mem[16710] = 'd0;
    mem[16711] = 'd512;
    mem[16712] = 'd0;
    mem[16713] = 'd872;
    mem[16714] = 'd0;
    mem[16715] = 'd0;
    mem[16716] = 'd0;
    mem[16717] = 'd524;
    mem[16718] = 'd0;
    mem[16719] = 'd876;
    mem[16720] = 'd0;
    mem[16721] = 'd0;
    mem[16722] = 'd0;
    mem[16723] = 'd528;
    mem[16724] = 'd0;
    mem[16725] = 'd880;
    mem[16726] = 'd0;
    mem[16727] = 'd0;
    mem[16728] = 'd0;
    mem[16729] = 'd528;
    mem[16730] = 'd0;
    mem[16731] = 'd880;
    mem[16732] = 'd0;
    mem[16733] = 'd0;
    mem[16734] = 'd0;
    mem[16735] = 'd524;
    mem[16736] = 'd0;
    mem[16737] = 'd876;
    mem[16738] = 'd0;
    mem[16739] = 'd0;
    mem[16740] = 'd0;
    mem[16741] = 'd512;
    mem[16742] = 'd0;
    mem[16743] = 'd872;
    mem[16744] = 'd0;
    mem[16745] = 'd0;
    mem[16746] = 'd0;
    mem[16747] = 'd496;
    mem[16748] = 'd0;
    mem[16749] = 'd860;
    mem[16750] = 'd0;
    mem[16751] = 'd0;
    mem[16752] = 'd0;
    mem[16753] = 'd472;
    mem[16754] = 'd0;
    mem[16755] = 'd840;
    mem[16756] = 'd0;
    mem[16757] = 'd0;
    mem[16758] = 'd0;
    mem[16759] = 'd436;
    mem[16760] = 'd0;
    mem[16761] = 'd804;
    mem[16762] = 'd0;
    mem[16763] = 'd0;
    mem[16764] = 'd0;
    mem[16765] = 'd608;
    mem[16766] = 'd0;
    mem[16767] = 'd860;
    mem[16768] = 'd0;
    mem[16769] = 'd0;
    mem[16770] = 'd0;
    mem[16771] = 'd836;
    mem[16772] = 'd0;
    mem[16773] = 'd948;
    mem[16774] = 'd0;
    mem[16775] = 'd0;
    mem[16776] = 'd0;
    mem[16777] = 'd996;
    mem[16778] = 'd0;
    mem[16779] = 'd1012;
    mem[16780] = 'd0;
    mem[16781] = 'd0;
    mem[16782] = 'd0;
    mem[16783] = 'd1016;
    mem[16784] = 'd0;
    mem[16785] = 'd1020;
    mem[16786] = 'd0;
    mem[16787] = 'd0;
    mem[16788] = 'd0;
    mem[16789] = 'd1020;
    mem[16790] = 'd0;
    mem[16791] = 'd1020;
    mem[16792] = 'd0;
    mem[16793] = 'd0;
    mem[16794] = 'd0;
    mem[16795] = 'd1020;
    mem[16796] = 'd0;
    mem[16797] = 'd1020;
    mem[16798] = 'd0;
    mem[16799] = 'd0;
    mem[16800] = 'd0;
    mem[16801] = 'd1020;
    mem[16802] = 'd0;
    mem[16803] = 'd1020;
    mem[16804] = 'd0;
    mem[16805] = 'd0;
    mem[16806] = 'd0;
    mem[16807] = 'd1020;
    mem[16808] = 'd0;
    mem[16809] = 'd1020;
    mem[16810] = 'd0;
    mem[16811] = 'd0;
    mem[16812] = 'd0;
    mem[16813] = 'd1020;
    mem[16814] = 'd0;
    mem[16815] = 'd1020;
    mem[16816] = 'd0;
    mem[16817] = 'd0;
    mem[16818] = 'd0;
    mem[16819] = 'd1020;
    mem[16820] = 'd0;
    mem[16821] = 'd1020;
    mem[16822] = 'd0;
    mem[16823] = 'd0;
    mem[16824] = 'd0;
    mem[16825] = 'd1020;
    mem[16826] = 'd0;
    mem[16827] = 'd1020;
    mem[16828] = 'd0;
    mem[16829] = 'd0;
    mem[16830] = 'd0;
    mem[16831] = 'd1020;
    mem[16832] = 'd0;
    mem[16833] = 'd1020;
    mem[16834] = 'd0;
    mem[16835] = 'd0;
    mem[16836] = 'd0;
    mem[16837] = 'd1020;
    mem[16838] = 'd0;
    mem[16839] = 'd1020;
    mem[16840] = 'd0;
    mem[16841] = 'd0;
    mem[16842] = 'd0;
    mem[16843] = 'd1020;
    mem[16844] = 'd0;
    mem[16845] = 'd1020;
    mem[16846] = 'd0;
    mem[16847] = 'd0;
    mem[16848] = 'd0;
    mem[16849] = 'd0;
    mem[16850] = 'd1020;
    mem[16851] = 'd0;
    mem[16852] = 'd1020;
    mem[16853] = 'd0;
    mem[16854] = 'd0;
    mem[16855] = 'd0;
    mem[16856] = 'd1020;
    mem[16857] = 'd0;
    mem[16858] = 'd1020;
    mem[16859] = 'd0;
    mem[16860] = 'd0;
    mem[16861] = 'd0;
    mem[16862] = 'd1020;
    mem[16863] = 'd0;
    mem[16864] = 'd1020;
    mem[16865] = 'd0;
    mem[16866] = 'd0;
    mem[16867] = 'd0;
    mem[16868] = 'd1020;
    mem[16869] = 'd0;
    mem[16870] = 'd1020;
    mem[16871] = 'd0;
    mem[16872] = 'd0;
    mem[16873] = 'd0;
    mem[16874] = 'd1020;
    mem[16875] = 'd0;
    mem[16876] = 'd1020;
    mem[16877] = 'd0;
    mem[16878] = 'd0;
    mem[16879] = 'd0;
    mem[16880] = 'd1020;
    mem[16881] = 'd0;
    mem[16882] = 'd1020;
    mem[16883] = 'd0;
    mem[16884] = 'd0;
    mem[16885] = 'd0;
    mem[16886] = 'd1020;
    mem[16887] = 'd0;
    mem[16888] = 'd1020;
    mem[16889] = 'd0;
    mem[16890] = 'd0;
    mem[16891] = 'd0;
    mem[16892] = 'd1020;
    mem[16893] = 'd0;
    mem[16894] = 'd1020;
    mem[16895] = 'd0;
    mem[16896] = 'd0;
    mem[16897] = 'd0;
    mem[16898] = 'd1020;
    mem[16899] = 'd0;
    mem[16900] = 'd1020;
    mem[16901] = 'd0;
    mem[16902] = 'd0;
    mem[16903] = 'd0;
    mem[16904] = 'd1016;
    mem[16905] = 'd0;
    mem[16906] = 'd1020;
    mem[16907] = 'd0;
    mem[16908] = 'd0;
    mem[16909] = 'd0;
    mem[16910] = 'd1012;
    mem[16911] = 'd0;
    mem[16912] = 'd1016;
    mem[16913] = 'd0;
    mem[16914] = 'd0;
    mem[16915] = 'd0;
    mem[16916] = 'd1012;
    mem[16917] = 'd0;
    mem[16918] = 'd1016;
    mem[16919] = 'd0;
    mem[16920] = 'd0;
    mem[16921] = 'd0;
    mem[16922] = 'd1008;
    mem[16923] = 'd0;
    mem[16924] = 'd1016;
    mem[16925] = 'd0;
    mem[16926] = 'd0;
    mem[16927] = 'd0;
    mem[16928] = 'd916;
    mem[16929] = 'd0;
    mem[16930] = 'd964;
    mem[16931] = 'd0;
    mem[16932] = 'd0;
    mem[16933] = 'd0;
    mem[16934] = 'd652;
    mem[16935] = 'd0;
    mem[16936] = 'd788;
    mem[16937] = 'd0;
    mem[16938] = 'd0;
    mem[16939] = 'd0;
    mem[16940] = 'd424;
    mem[16941] = 'd0;
    mem[16942] = 'd652;
    mem[16943] = 'd0;
    mem[16944] = 'd0;
    mem[16945] = 'd0;
    mem[16946] = 'd252;
    mem[16947] = 'd0;
    mem[16948] = 'd556;
    mem[16949] = 'd0;
    mem[16950] = 'd0;
    mem[16951] = 'd0;
    mem[16952] = 'd148;
    mem[16953] = 'd0;
    mem[16954] = 'd496;
    mem[16955] = 'd0;
    mem[16956] = 'd0;
    mem[16957] = 'd0;
    mem[16958] = 'd100;
    mem[16959] = 'd0;
    mem[16960] = 'd472;
    mem[16961] = 'd0;
    mem[16962] = 'd0;
    mem[16963] = 'd0;
    mem[16964] = 'd100;
    mem[16965] = 'd0;
    mem[16966] = 'd472;
    mem[16967] = 'd0;
    mem[16968] = 'd0;
    mem[16969] = 'd0;
    mem[16970] = 'd144;
    mem[16971] = 'd0;
    mem[16972] = 'd496;
    mem[16973] = 'd0;
    mem[16974] = 'd0;
    mem[16975] = 'd0;
    mem[16976] = 'd248;
    mem[16977] = 'd0;
    mem[16978] = 'd552;
    mem[16979] = 'd0;
    mem[16980] = 'd0;
    mem[16981] = 'd0;
    mem[16982] = 'd416;
    mem[16983] = 'd0;
    mem[16984] = 'd648;
    mem[16985] = 'd0;
    mem[16986] = 'd0;
    mem[16987] = 'd0;
    mem[16988] = 'd652;
    mem[16989] = 'd0;
    mem[16990] = 'd792;
    mem[16991] = 'd0;
    mem[16992] = 'd0;
    mem[16993] = 'd0;
    mem[16994] = 'd952;
    mem[16995] = 'd0;
    mem[16996] = 'd984;
    mem[16997] = 'd0;
    mem[16998] = 'd0;
    mem[16999] = 'd0;
    mem[17000] = 'd1004;
    mem[17001] = 'd0;
    mem[17002] = 'd1016;
    mem[17003] = 'd0;
    mem[17004] = 'd0;
    mem[17005] = 'd0;
    mem[17006] = 'd1012;
    mem[17007] = 'd0;
    mem[17008] = 'd1016;
    mem[17009] = 'd0;
    mem[17010] = 'd0;
    mem[17011] = 'd0;
    mem[17012] = 'd1016;
    mem[17013] = 'd0;
    mem[17014] = 'd1020;
    mem[17015] = 'd0;
    mem[17016] = 'd0;
    mem[17017] = 'd0;
    mem[17018] = 'd1016;
    mem[17019] = 'd0;
    mem[17020] = 'd1020;
    mem[17021] = 'd0;
    mem[17022] = 'd0;
    mem[17023] = 'd0;
    mem[17024] = 'd1020;
    mem[17025] = 'd0;
    mem[17026] = 'd1020;
    mem[17027] = 'd0;
    mem[17028] = 'd0;
    mem[17029] = 'd0;
    mem[17030] = 'd1020;
    mem[17031] = 'd0;
    mem[17032] = 'd1020;
    mem[17033] = 'd0;
    mem[17034] = 'd0;
    mem[17035] = 'd0;
    mem[17036] = 'd1020;
    mem[17037] = 'd0;
    mem[17038] = 'd1020;
    mem[17039] = 'd0;
    mem[17040] = 'd0;
    mem[17041] = 'd0;
    mem[17042] = 'd1020;
    mem[17043] = 'd0;
    mem[17044] = 'd1020;
    mem[17045] = 'd0;
    mem[17046] = 'd0;
    mem[17047] = 'd0;
    mem[17048] = 'd1020;
    mem[17049] = 'd0;
    mem[17050] = 'd1020;
    mem[17051] = 'd0;
    mem[17052] = 'd0;
    mem[17053] = 'd0;
    mem[17054] = 'd1020;
    mem[17055] = 'd0;
    mem[17056] = 'd1020;
    mem[17057] = 'd0;
    mem[17058] = 'd0;
    mem[17059] = 'd0;
    mem[17060] = 'd1020;
    mem[17061] = 'd0;
    mem[17062] = 'd1020;
    mem[17063] = 'd0;
    mem[17064] = 'd0;
    mem[17065] = 'd0;
    mem[17066] = 'd1020;
    mem[17067] = 'd0;
    mem[17068] = 'd1020;
    mem[17069] = 'd0;
    mem[17070] = 'd0;
    mem[17071] = 'd0;
    mem[17072] = 'd1020;
    mem[17073] = 'd0;
    mem[17074] = 'd1020;
    mem[17075] = 'd0;
    mem[17076] = 'd0;
    mem[17077] = 'd0;
    mem[17078] = 'd1020;
    mem[17079] = 'd0;
    mem[17080] = 'd1020;
    mem[17081] = 'd0;
    mem[17082] = 'd0;
    mem[17083] = 'd1020;
    mem[17084] = 'd0;
    mem[17085] = 'd1020;
    mem[17086] = 'd0;
    mem[17087] = 'd0;
    mem[17088] = 'd0;
    mem[17089] = 'd1020;
    mem[17090] = 'd0;
    mem[17091] = 'd1020;
    mem[17092] = 'd0;
    mem[17093] = 'd0;
    mem[17094] = 'd0;
    mem[17095] = 'd1020;
    mem[17096] = 'd0;
    mem[17097] = 'd1020;
    mem[17098] = 'd0;
    mem[17099] = 'd0;
    mem[17100] = 'd0;
    mem[17101] = 'd1020;
    mem[17102] = 'd0;
    mem[17103] = 'd1020;
    mem[17104] = 'd0;
    mem[17105] = 'd0;
    mem[17106] = 'd0;
    mem[17107] = 'd1020;
    mem[17108] = 'd0;
    mem[17109] = 'd1020;
    mem[17110] = 'd0;
    mem[17111] = 'd0;
    mem[17112] = 'd0;
    mem[17113] = 'd1020;
    mem[17114] = 'd0;
    mem[17115] = 'd1020;
    mem[17116] = 'd0;
    mem[17117] = 'd0;
    mem[17118] = 'd0;
    mem[17119] = 'd1020;
    mem[17120] = 'd0;
    mem[17121] = 'd1020;
    mem[17122] = 'd0;
    mem[17123] = 'd0;
    mem[17124] = 'd0;
    mem[17125] = 'd1020;
    mem[17126] = 'd0;
    mem[17127] = 'd1020;
    mem[17128] = 'd0;
    mem[17129] = 'd0;
    mem[17130] = 'd0;
    mem[17131] = 'd1020;
    mem[17132] = 'd0;
    mem[17133] = 'd1020;
    mem[17134] = 'd0;
    mem[17135] = 'd0;
    mem[17136] = 'd0;
    mem[17137] = 'd1020;
    mem[17138] = 'd0;
    mem[17139] = 'd1020;
    mem[17140] = 'd0;
    mem[17141] = 'd0;
    mem[17142] = 'd0;
    mem[17143] = 'd1016;
    mem[17144] = 'd0;
    mem[17145] = 'd1020;
    mem[17146] = 'd0;
    mem[17147] = 'd0;
    mem[17148] = 'd0;
    mem[17149] = 'd1016;
    mem[17150] = 'd0;
    mem[17151] = 'd1020;
    mem[17152] = 'd0;
    mem[17153] = 'd0;
    mem[17154] = 'd0;
    mem[17155] = 'd1016;
    mem[17156] = 'd0;
    mem[17157] = 'd1020;
    mem[17158] = 'd0;
    mem[17159] = 'd0;
    mem[17160] = 'd0;
    mem[17161] = 'd964;
    mem[17162] = 'd0;
    mem[17163] = 'd996;
    mem[17164] = 'd0;
    mem[17165] = 'd0;
    mem[17166] = 'd0;
    mem[17167] = 'd788;
    mem[17168] = 'd0;
    mem[17169] = 'd924;
    mem[17170] = 'd0;
    mem[17171] = 'd0;
    mem[17172] = 'd0;
    mem[17173] = 'd652;
    mem[17174] = 'd0;
    mem[17175] = 'd868;
    mem[17176] = 'd0;
    mem[17177] = 'd0;
    mem[17178] = 'd0;
    mem[17179] = 'd556;
    mem[17180] = 'd0;
    mem[17181] = 'd836;
    mem[17182] = 'd0;
    mem[17183] = 'd0;
    mem[17184] = 'd0;
    mem[17185] = 'd496;
    mem[17186] = 'd0;
    mem[17187] = 'd816;
    mem[17188] = 'd0;
    mem[17189] = 'd0;
    mem[17190] = 'd0;
    mem[17191] = 'd472;
    mem[17192] = 'd0;
    mem[17193] = 'd808;
    mem[17194] = 'd0;
    mem[17195] = 'd0;
    mem[17196] = 'd0;
    mem[17197] = 'd472;
    mem[17198] = 'd0;
    mem[17199] = 'd808;
    mem[17200] = 'd0;
    mem[17201] = 'd0;
    mem[17202] = 'd0;
    mem[17203] = 'd496;
    mem[17204] = 'd0;
    mem[17205] = 'd816;
    mem[17206] = 'd0;
    mem[17207] = 'd0;
    mem[17208] = 'd0;
    mem[17209] = 'd552;
    mem[17210] = 'd0;
    mem[17211] = 'd836;
    mem[17212] = 'd0;
    mem[17213] = 'd0;
    mem[17214] = 'd0;
    mem[17215] = 'd648;
    mem[17216] = 'd0;
    mem[17217] = 'd868;
    mem[17218] = 'd0;
    mem[17219] = 'd0;
    mem[17220] = 'd0;
    mem[17221] = 'd792;
    mem[17222] = 'd0;
    mem[17223] = 'd920;
    mem[17224] = 'd0;
    mem[17225] = 'd0;
    mem[17226] = 'd0;
    mem[17227] = 'd984;
    mem[17228] = 'd0;
    mem[17229] = 'd1008;
    mem[17230] = 'd0;
    mem[17231] = 'd0;
    mem[17232] = 'd0;
    mem[17233] = 'd1016;
    mem[17234] = 'd0;
    mem[17235] = 'd1020;
    mem[17236] = 'd0;
    mem[17237] = 'd0;
    mem[17238] = 'd0;
    mem[17239] = 'd1016;
    mem[17240] = 'd0;
    mem[17241] = 'd1020;
    mem[17242] = 'd0;
    mem[17243] = 'd0;
    mem[17244] = 'd0;
    mem[17245] = 'd1020;
    mem[17246] = 'd0;
    mem[17247] = 'd1020;
    mem[17248] = 'd0;
    mem[17249] = 'd0;
    mem[17250] = 'd0;
    mem[17251] = 'd1020;
    mem[17252] = 'd0;
    mem[17253] = 'd1020;
    mem[17254] = 'd0;
    mem[17255] = 'd0;
    mem[17256] = 'd0;
    mem[17257] = 'd1020;
    mem[17258] = 'd0;
    mem[17259] = 'd1020;
    mem[17260] = 'd0;
    mem[17261] = 'd0;
    mem[17262] = 'd0;
    mem[17263] = 'd1020;
    mem[17264] = 'd0;
    mem[17265] = 'd1020;
    mem[17266] = 'd0;
    mem[17267] = 'd0;
    mem[17268] = 'd0;
    mem[17269] = 'd1020;
    mem[17270] = 'd0;
    mem[17271] = 'd1020;
    mem[17272] = 'd0;
    mem[17273] = 'd0;
    mem[17274] = 'd0;
    mem[17275] = 'd1020;
    mem[17276] = 'd0;
    mem[17277] = 'd1020;
    mem[17278] = 'd0;
    mem[17279] = 'd0;
    mem[17280] = 'd0;
    mem[17281] = 'd1020;
    mem[17282] = 'd0;
    mem[17283] = 'd1020;
    mem[17284] = 'd0;
    mem[17285] = 'd0;
    mem[17286] = 'd0;
    mem[17287] = 'd1020;
    mem[17288] = 'd0;
    mem[17289] = 'd1020;
    mem[17290] = 'd0;
    mem[17291] = 'd0;
    mem[17292] = 'd0;
    mem[17293] = 'd1020;
    mem[17294] = 'd0;
    mem[17295] = 'd1020;
    mem[17296] = 'd0;
    mem[17297] = 'd0;
    mem[17298] = 'd0;
    mem[17299] = 'd1020;
    mem[17300] = 'd0;
    mem[17301] = 'd1020;
    mem[17302] = 'd0;
    mem[17303] = 'd0;
    mem[17304] = 'd0;
    mem[17305] = 'd1020;
    mem[17306] = 'd0;
    mem[17307] = 'd1020;
    mem[17308] = 'd0;
    mem[17309] = 'd0;
    mem[17310] = 'd0;
    mem[17311] = 'd1020;
    mem[17312] = 'd0;
    mem[17313] = 'd1020;
    mem[17314] = 'd0;
    mem[17315] = 'd0;
    mem[17316] = 'd0;
    mem[17317] = 'd0;
    mem[17318] = 'd1020;
    mem[17319] = 'd0;
    mem[17320] = 'd1020;
    mem[17321] = 'd0;
    mem[17322] = 'd0;
    mem[17323] = 'd0;
    mem[17324] = 'd1020;
    mem[17325] = 'd0;
    mem[17326] = 'd1020;
    mem[17327] = 'd0;
    mem[17328] = 'd0;
    mem[17329] = 'd0;
    mem[17330] = 'd1020;
    mem[17331] = 'd0;
    mem[17332] = 'd1020;
    mem[17333] = 'd0;
    mem[17334] = 'd0;
    mem[17335] = 'd0;
    mem[17336] = 'd1020;
    mem[17337] = 'd0;
    mem[17338] = 'd1020;
    mem[17339] = 'd0;
    mem[17340] = 'd0;
    mem[17341] = 'd0;
    mem[17342] = 'd1020;
    mem[17343] = 'd0;
    mem[17344] = 'd1020;
    mem[17345] = 'd0;
    mem[17346] = 'd0;
    mem[17347] = 'd0;
    mem[17348] = 'd1020;
    mem[17349] = 'd0;
    mem[17350] = 'd1020;
    mem[17351] = 'd0;
    mem[17352] = 'd0;
    mem[17353] = 'd0;
    mem[17354] = 'd1020;
    mem[17355] = 'd0;
    mem[17356] = 'd1020;
    mem[17357] = 'd0;
    mem[17358] = 'd0;
    mem[17359] = 'd0;
    mem[17360] = 'd1020;
    mem[17361] = 'd0;
    mem[17362] = 'd1020;
    mem[17363] = 'd0;
    mem[17364] = 'd0;
    mem[17365] = 'd0;
    mem[17366] = 'd1020;
    mem[17367] = 'd0;
    mem[17368] = 'd1020;
    mem[17369] = 'd0;
    mem[17370] = 'd0;
    mem[17371] = 'd0;
    mem[17372] = 'd1020;
    mem[17373] = 'd0;
    mem[17374] = 'd1020;
    mem[17375] = 'd0;
    mem[17376] = 'd0;
    mem[17377] = 'd0;
    mem[17378] = 'd1020;
    mem[17379] = 'd0;
    mem[17380] = 'd1020;
    mem[17381] = 'd0;
    mem[17382] = 'd0;
    mem[17383] = 'd0;
    mem[17384] = 'd1016;
    mem[17385] = 'd0;
    mem[17386] = 'd1020;
    mem[17387] = 'd0;
    mem[17388] = 'd0;
    mem[17389] = 'd0;
    mem[17390] = 'd1016;
    mem[17391] = 'd0;
    mem[17392] = 'd1020;
    mem[17393] = 'd0;
    mem[17394] = 'd0;
    mem[17395] = 'd0;
    mem[17396] = 'd1012;
    mem[17397] = 'd0;
    mem[17398] = 'd1016;
    mem[17399] = 'd0;
    mem[17400] = 'd0;
    mem[17401] = 'd0;
    mem[17402] = 'd1012;
    mem[17403] = 'd0;
    mem[17404] = 'd1016;
    mem[17405] = 'd0;
    mem[17406] = 'd0;
    mem[17407] = 'd0;
    mem[17408] = 'd1008;
    mem[17409] = 'd0;
    mem[17410] = 'd1016;
    mem[17411] = 'd0;
    mem[17412] = 'd0;
    mem[17413] = 'd0;
    mem[17414] = 'd1008;
    mem[17415] = 'd0;
    mem[17416] = 'd1016;
    mem[17417] = 'd0;
    mem[17418] = 'd0;
    mem[17419] = 'd0;
    mem[17420] = 'd1008;
    mem[17421] = 'd0;
    mem[17422] = 'd1016;
    mem[17423] = 'd0;
    mem[17424] = 'd0;
    mem[17425] = 'd0;
    mem[17426] = 'd1004;
    mem[17427] = 'd0;
    mem[17428] = 'd1012;
    mem[17429] = 'd0;
    mem[17430] = 'd0;
    mem[17431] = 'd0;
    mem[17432] = 'd1000;
    mem[17433] = 'd0;
    mem[17434] = 'd1012;
    mem[17435] = 'd0;
    mem[17436] = 'd0;
    mem[17437] = 'd0;
    mem[17438] = 'd1008;
    mem[17439] = 'd0;
    mem[17440] = 'd1016;
    mem[17441] = 'd0;
    mem[17442] = 'd0;
    mem[17443] = 'd0;
    mem[17444] = 'd1008;
    mem[17445] = 'd0;
    mem[17446] = 'd1016;
    mem[17447] = 'd0;
    mem[17448] = 'd0;
    mem[17449] = 'd0;
    mem[17450] = 'd1008;
    mem[17451] = 'd0;
    mem[17452] = 'd1016;
    mem[17453] = 'd0;
    mem[17454] = 'd0;
    mem[17455] = 'd0;
    mem[17456] = 'd1008;
    mem[17457] = 'd0;
    mem[17458] = 'd1016;
    mem[17459] = 'd0;
    mem[17460] = 'd0;
    mem[17461] = 'd0;
    mem[17462] = 'd1012;
    mem[17463] = 'd0;
    mem[17464] = 'd1016;
    mem[17465] = 'd0;
    mem[17466] = 'd0;
    mem[17467] = 'd0;
    mem[17468] = 'd1016;
    mem[17469] = 'd0;
    mem[17470] = 'd1020;
    mem[17471] = 'd0;
    mem[17472] = 'd0;
    mem[17473] = 'd0;
    mem[17474] = 'd1016;
    mem[17475] = 'd0;
    mem[17476] = 'd1020;
    mem[17477] = 'd0;
    mem[17478] = 'd0;
    mem[17479] = 'd0;
    mem[17480] = 'd1020;
    mem[17481] = 'd0;
    mem[17482] = 'd1020;
    mem[17483] = 'd0;
    mem[17484] = 'd0;
    mem[17485] = 'd0;
    mem[17486] = 'd1020;
    mem[17487] = 'd0;
    mem[17488] = 'd1020;
    mem[17489] = 'd0;
    mem[17490] = 'd0;
    mem[17491] = 'd0;
    mem[17492] = 'd1020;
    mem[17493] = 'd0;
    mem[17494] = 'd1020;
    mem[17495] = 'd0;
    mem[17496] = 'd0;
    mem[17497] = 'd0;
    mem[17498] = 'd1020;
    mem[17499] = 'd0;
    mem[17500] = 'd1020;
    mem[17501] = 'd0;
    mem[17502] = 'd0;
    mem[17503] = 'd0;
    mem[17504] = 'd1020;
    mem[17505] = 'd0;
    mem[17506] = 'd1020;
    mem[17507] = 'd0;
    mem[17508] = 'd0;
    mem[17509] = 'd0;
    mem[17510] = 'd1020;
    mem[17511] = 'd0;
    mem[17512] = 'd1020;
    mem[17513] = 'd0;
    mem[17514] = 'd0;
    mem[17515] = 'd0;
    mem[17516] = 'd1020;
    mem[17517] = 'd0;
    mem[17518] = 'd1020;
    mem[17519] = 'd0;
    mem[17520] = 'd0;
    mem[17521] = 'd0;
    mem[17522] = 'd1020;
    mem[17523] = 'd0;
    mem[17524] = 'd1020;
    mem[17525] = 'd0;
    mem[17526] = 'd0;
    mem[17527] = 'd0;
    mem[17528] = 'd1020;
    mem[17529] = 'd0;
    mem[17530] = 'd1020;
    mem[17531] = 'd0;
    mem[17532] = 'd0;
    mem[17533] = 'd0;
    mem[17534] = 'd1020;
    mem[17535] = 'd0;
    mem[17536] = 'd1020;
    mem[17537] = 'd0;
    mem[17538] = 'd0;
    mem[17539] = 'd0;
    mem[17540] = 'd1020;
    mem[17541] = 'd0;
    mem[17542] = 'd1020;
    mem[17543] = 'd0;
    mem[17544] = 'd0;
    mem[17545] = 'd0;
    mem[17546] = 'd1020;
    mem[17547] = 'd0;
    mem[17548] = 'd1020;
    mem[17549] = 'd0;
    mem[17550] = 'd0;
    mem[17551] = 'd1020;
    mem[17552] = 'd0;
    mem[17553] = 'd1020;
    mem[17554] = 'd0;
    mem[17555] = 'd0;
    mem[17556] = 'd0;
    mem[17557] = 'd1020;
    mem[17558] = 'd0;
    mem[17559] = 'd1020;
    mem[17560] = 'd0;
    mem[17561] = 'd0;
    mem[17562] = 'd0;
    mem[17563] = 'd1020;
    mem[17564] = 'd0;
    mem[17565] = 'd1020;
    mem[17566] = 'd0;
    mem[17567] = 'd0;
    mem[17568] = 'd0;
    mem[17569] = 'd1020;
    mem[17570] = 'd0;
    mem[17571] = 'd1020;
    mem[17572] = 'd0;
    mem[17573] = 'd0;
    mem[17574] = 'd0;
    mem[17575] = 'd1020;
    mem[17576] = 'd0;
    mem[17577] = 'd1020;
    mem[17578] = 'd0;
    mem[17579] = 'd0;
    mem[17580] = 'd0;
    mem[17581] = 'd1020;
    mem[17582] = 'd0;
    mem[17583] = 'd1020;
    mem[17584] = 'd0;
    mem[17585] = 'd0;
    mem[17586] = 'd0;
    mem[17587] = 'd1020;
    mem[17588] = 'd0;
    mem[17589] = 'd1020;
    mem[17590] = 'd0;
    mem[17591] = 'd0;
    mem[17592] = 'd0;
    mem[17593] = 'd1020;
    mem[17594] = 'd0;
    mem[17595] = 'd1020;
    mem[17596] = 'd0;
    mem[17597] = 'd0;
    mem[17598] = 'd0;
    mem[17599] = 'd1020;
    mem[17600] = 'd0;
    mem[17601] = 'd1020;
    mem[17602] = 'd0;
    mem[17603] = 'd0;
    mem[17604] = 'd0;
    mem[17605] = 'd1020;
    mem[17606] = 'd0;
    mem[17607] = 'd1020;
    mem[17608] = 'd0;
    mem[17609] = 'd0;
    mem[17610] = 'd0;
    mem[17611] = 'd1020;
    mem[17612] = 'd0;
    mem[17613] = 'd1020;
    mem[17614] = 'd0;
    mem[17615] = 'd0;
    mem[17616] = 'd0;
    mem[17617] = 'd1020;
    mem[17618] = 'd0;
    mem[17619] = 'd1020;
    mem[17620] = 'd0;
    mem[17621] = 'd0;
    mem[17622] = 'd0;
    mem[17623] = 'd1020;
    mem[17624] = 'd0;
    mem[17625] = 'd1020;
    mem[17626] = 'd0;
    mem[17627] = 'd0;
    mem[17628] = 'd0;
    mem[17629] = 'd1016;
    mem[17630] = 'd0;
    mem[17631] = 'd1020;
    mem[17632] = 'd0;
    mem[17633] = 'd0;
    mem[17634] = 'd0;
    mem[17635] = 'd1016;
    mem[17636] = 'd0;
    mem[17637] = 'd1020;
    mem[17638] = 'd0;
    mem[17639] = 'd0;
    mem[17640] = 'd0;
    mem[17641] = 'd1016;
    mem[17642] = 'd0;
    mem[17643] = 'd1020;
    mem[17644] = 'd0;
    mem[17645] = 'd0;
    mem[17646] = 'd0;
    mem[17647] = 'd1016;
    mem[17648] = 'd0;
    mem[17649] = 'd1020;
    mem[17650] = 'd0;
    mem[17651] = 'd0;
    mem[17652] = 'd0;
    mem[17653] = 'd1016;
    mem[17654] = 'd0;
    mem[17655] = 'd1020;
    mem[17656] = 'd0;
    mem[17657] = 'd0;
    mem[17658] = 'd0;
    mem[17659] = 'd1012;
    mem[17660] = 'd0;
    mem[17661] = 'd1020;
    mem[17662] = 'd0;
    mem[17663] = 'd0;
    mem[17664] = 'd0;
    mem[17665] = 'd1012;
    mem[17666] = 'd0;
    mem[17667] = 'd1020;
    mem[17668] = 'd0;
    mem[17669] = 'd0;
    mem[17670] = 'd0;
    mem[17671] = 'd1016;
    mem[17672] = 'd0;
    mem[17673] = 'd1020;
    mem[17674] = 'd0;
    mem[17675] = 'd0;
    mem[17676] = 'd0;
    mem[17677] = 'd1016;
    mem[17678] = 'd0;
    mem[17679] = 'd1020;
    mem[17680] = 'd0;
    mem[17681] = 'd0;
    mem[17682] = 'd0;
    mem[17683] = 'd1016;
    mem[17684] = 'd0;
    mem[17685] = 'd1020;
    mem[17686] = 'd0;
    mem[17687] = 'd0;
    mem[17688] = 'd0;
    mem[17689] = 'd1016;
    mem[17690] = 'd0;
    mem[17691] = 'd1020;
    mem[17692] = 'd0;
    mem[17693] = 'd0;
    mem[17694] = 'd0;
    mem[17695] = 'd1016;
    mem[17696] = 'd0;
    mem[17697] = 'd1020;
    mem[17698] = 'd0;
    mem[17699] = 'd0;
    mem[17700] = 'd0;
    mem[17701] = 'd1020;
    mem[17702] = 'd0;
    mem[17703] = 'd1020;
    mem[17704] = 'd0;
    mem[17705] = 'd0;
    mem[17706] = 'd0;
    mem[17707] = 'd1020;
    mem[17708] = 'd0;
    mem[17709] = 'd1020;
    mem[17710] = 'd0;
    mem[17711] = 'd0;
    mem[17712] = 'd0;
    mem[17713] = 'd1020;
    mem[17714] = 'd0;
    mem[17715] = 'd1020;
    mem[17716] = 'd0;
    mem[17717] = 'd0;
    mem[17718] = 'd0;
    mem[17719] = 'd1020;
    mem[17720] = 'd0;
    mem[17721] = 'd1020;
    mem[17722] = 'd0;
    mem[17723] = 'd0;
    mem[17724] = 'd0;
    mem[17725] = 'd1020;
    mem[17726] = 'd0;
    mem[17727] = 'd1020;
    mem[17728] = 'd0;
    mem[17729] = 'd0;
    mem[17730] = 'd0;
    mem[17731] = 'd1020;
    mem[17732] = 'd0;
    mem[17733] = 'd1020;
    mem[17734] = 'd0;
    mem[17735] = 'd0;
    mem[17736] = 'd0;
    mem[17737] = 'd1020;
    mem[17738] = 'd0;
    mem[17739] = 'd1020;
    mem[17740] = 'd0;
    mem[17741] = 'd0;
    mem[17742] = 'd0;
    mem[17743] = 'd1020;
    mem[17744] = 'd0;
    mem[17745] = 'd1020;
    mem[17746] = 'd0;
    mem[17747] = 'd0;
    mem[17748] = 'd0;
    mem[17749] = 'd1020;
    mem[17750] = 'd0;
    mem[17751] = 'd1020;
    mem[17752] = 'd0;
    mem[17753] = 'd0;
    mem[17754] = 'd0;
    mem[17755] = 'd1020;
    mem[17756] = 'd0;
    mem[17757] = 'd1020;
    mem[17758] = 'd0;
    mem[17759] = 'd0;
    mem[17760] = 'd0;
    mem[17761] = 'd1020;
    mem[17762] = 'd0;
    mem[17763] = 'd1020;
    mem[17764] = 'd0;
    mem[17765] = 'd0;
    mem[17766] = 'd0;
    mem[17767] = 'd1020;
    mem[17768] = 'd0;
    mem[17769] = 'd1020;
    mem[17770] = 'd0;
    mem[17771] = 'd0;
    mem[17772] = 'd0;
    mem[17773] = 'd1020;
    mem[17774] = 'd0;
    mem[17775] = 'd1020;
    mem[17776] = 'd0;
    mem[17777] = 'd0;
    mem[17778] = 'd0;
    mem[17779] = 'd1020;
    mem[17780] = 'd0;
    mem[17781] = 'd1020;
    mem[17782] = 'd0;
    mem[17783] = 'd0;

end

endmodule