/*
 * This file is a part of: https://github.com/brilliantlabsAR/frame-codebase
 *
 * Authored by: Rohit Rathnam / Silicon Witchery AB (rohit@siliconwitchery.com)
 *              Raj Nakarja / Brilliant Labs Limited (raj@brilliant.xyz)
 *
 * CERN Open Hardware Licence Version 2 - Permissive
 *
 * Copyright © 2023 Brilliant Labs Limited
 */

module image_gen #(
    parameter X_RESOLUTION = 78,
    parameter Y_RESOLUTION = 76,
    parameter H_FRONT_PORCH = 156, // 2x X_RESOLUTION
    parameter H_BACK_PORCH = 172, // ~ 2.2x X_RESOLUTION
    parameter V_FRONT_PORCH = 1,
    parameter V_BACK_PORCH = 2,
    parameter H_SYNC_PULSE_WIDTH = 44,
    parameter V_SYNC_PULSE_WIDTH = 5
) (
    input logic pixel_clock_in,
    input logic reset_n_in,

    output logic [9:0] pixel_data_out,
    output logic line_valid,
    output logic frame_valid
);

logic [31:0] x_counter;
logic [31:0] y_counter;
logic [31:0] pixel_counter;

logic [9:0] mem[5927:0];

always @(posedge pixel_clock_in) begin

    if(!reset_n_in) begin

        pixel_data_out <= 0;
        line_valid <= 0;
        frame_valid <= 0;

        x_counter <= 0;
        y_counter <= 0;
        pixel_counter <= 0;

    end 

    else begin
            
        // Increment counters
        if (x_counter <= (H_SYNC_PULSE_WIDTH + H_BACK_PORCH + X_RESOLUTION + H_FRONT_PORCH)) begin
            x_counter <= x_counter + 1;
        end

        else begin
            x_counter <= 0;

            if (y_counter <= (V_SYNC_PULSE_WIDTH + V_BACK_PORCH + Y_RESOLUTION + V_FRONT_PORCH)) begin
                y_counter <= y_counter + 1;
            end

            else begin
                y_counter <= 0;
            end 

        end

        // Output line valud
        if ((x_counter >= (H_SYNC_PULSE_WIDTH + H_BACK_PORCH)) &&
            (x_counter < (H_SYNC_PULSE_WIDTH + H_BACK_PORCH + X_RESOLUTION)) &&
            (y_counter >= (V_SYNC_PULSE_WIDTH + V_BACK_PORCH)) &&
            (y_counter < (V_SYNC_PULSE_WIDTH + V_BACK_PORCH + Y_RESOLUTION))) begin
                
            line_valid <= 1;

            pixel_counter <= pixel_counter + 1;
        end

        else begin
            line_valid <= 0;
        end

        // Output frame valid
        if (y_counter >= 0 &&
            y_counter < V_SYNC_PULSE_WIDTH) begin

            frame_valid <= 0;
            pixel_counter <= 0;

        end

        else begin
            frame_valid <= 1;
        end
        
        // Output pixel
        pixel_data_out <= mem[pixel_counter];

    end

end

initial begin

    mem[0] = 'd1020;
    mem[1] = 'd1020;
    mem[2] = 'd1020;
    mem[3] = 'd1020;
    mem[4] = 'd1020;
    mem[5] = 'd1020;
    mem[6] = 'd1020;
    mem[7] = 'd1020;
    mem[8] = 'd1020;
    mem[9] = 'd1020;
    mem[10] = 'd1020;
    mem[11] = 'd1020;
    mem[12] = 'd1020;
    mem[13] = 'd1020;
    mem[14] = 'd1020;
    mem[15] = 'd1020;
    mem[16] = 'd1020;
    mem[17] = 'd1020;
    mem[18] = 'd1020;
    mem[19] = 'd1020;
    mem[20] = 'd1020;
    mem[21] = 'd1020;
    mem[22] = 'd1020;
    mem[23] = 'd1020;
    mem[24] = 'd1020;
    mem[25] = 'd1020;
    mem[26] = 'd1020;
    mem[27] = 'd1020;
    mem[28] = 'd1020;
    mem[29] = 'd1020;
    mem[30] = 'd1020;
    mem[31] = 'd1020;
    mem[32] = 'd1020;
    mem[33] = 'd1020;
    mem[34] = 'd1020;
    mem[35] = 'd1020;
    mem[36] = 'd1020;
    mem[37] = 'd1020;
    mem[38] = 'd1020;
    mem[39] = 'd1020;
    mem[40] = 'd1020;
    mem[41] = 'd1020;
    mem[42] = 'd1020;
    mem[43] = 'd1020;
    mem[44] = 'd1020;
    mem[45] = 'd1020;
    mem[46] = 'd1020;
    mem[47] = 'd1020;
    mem[48] = 'd1020;
    mem[49] = 'd1020;
    mem[50] = 'd1020;
    mem[51] = 'd1020;
    mem[52] = 'd1020;
    mem[53] = 'd1020;
    mem[54] = 'd1020;
    mem[55] = 'd1020;
    mem[56] = 'd1020;
    mem[57] = 'd1020;
    mem[58] = 'd1020;
    mem[59] = 'd1020;
    mem[60] = 'd1020;
    mem[61] = 'd1020;
    mem[62] = 'd1020;
    mem[63] = 'd1020;
    mem[64] = 'd1020;
    mem[65] = 'd1020;
    mem[66] = 'd1020;
    mem[67] = 'd1020;
    mem[68] = 'd1020;
    mem[69] = 'd1020;
    mem[70] = 'd1020;
    mem[71] = 'd1020;
    mem[72] = 'd1020;
    mem[73] = 'd1020;
    mem[74] = 'd1020;
    mem[75] = 'd1020;
    mem[76] = 'd1020;
    mem[77] = 'd1020;
    mem[78] = 'd1020;
    mem[79] = 'd1020;
    mem[80] = 'd1020;
    mem[81] = 'd1020;
    mem[82] = 'd1020;
    mem[83] = 'd1020;
    mem[84] = 'd1020;
    mem[85] = 'd1020;
    mem[86] = 'd1020;
    mem[87] = 'd1020;
    mem[88] = 'd1020;
    mem[89] = 'd1020;
    mem[90] = 'd1020;
    mem[91] = 'd1020;
    mem[92] = 'd1020;
    mem[93] = 'd1020;
    mem[94] = 'd1020;
    mem[95] = 'd1020;
    mem[96] = 'd1020;
    mem[97] = 'd1020;
    mem[98] = 'd1020;
    mem[99] = 'd1020;
    mem[100] = 'd1020;
    mem[101] = 'd1020;
    mem[102] = 'd1020;
    mem[103] = 'd1020;
    mem[104] = 'd1020;
    mem[105] = 'd1020;
    mem[106] = 'd1020;
    mem[107] = 'd1020;
    mem[108] = 'd1020;
    mem[109] = 'd1020;
    mem[110] = 'd1020;
    mem[111] = 'd1020;
    mem[112] = 'd1020;
    mem[113] = 'd1020;
    mem[114] = 'd1020;
    mem[115] = 'd1020;
    mem[116] = 'd1020;
    mem[117] = 'd1020;
    mem[118] = 'd1020;
    mem[119] = 'd1020;
    mem[120] = 'd1020;
    mem[121] = 'd1020;
    mem[122] = 'd1020;
    mem[123] = 'd1020;
    mem[124] = 'd1020;
    mem[125] = 'd1020;
    mem[126] = 'd1020;
    mem[127] = 'd1020;
    mem[128] = 'd1020;
    mem[129] = 'd1020;
    mem[130] = 'd1020;
    mem[131] = 'd1020;
    mem[132] = 'd1020;
    mem[133] = 'd1020;
    mem[134] = 'd1020;
    mem[135] = 'd1020;
    mem[136] = 'd1020;
    mem[137] = 'd1020;
    mem[138] = 'd1020;
    mem[139] = 'd1020;
    mem[140] = 'd1020;
    mem[141] = 'd1020;
    mem[142] = 'd1020;
    mem[143] = 'd1020;
    mem[144] = 'd1020;
    mem[145] = 'd1020;
    mem[146] = 'd1020;
    mem[147] = 'd1020;
    mem[148] = 'd1020;
    mem[149] = 'd1020;
    mem[150] = 'd1020;
    mem[151] = 'd1020;
    mem[152] = 'd1020;
    mem[153] = 'd1020;
    mem[154] = 'd1020;
    mem[155] = 'd1020;
    mem[156] = 'd1020;
    mem[157] = 'd1020;
    mem[158] = 'd1020;
    mem[159] = 'd1020;
    mem[160] = 'd1020;
    mem[161] = 'd1020;
    mem[162] = 'd1020;
    mem[163] = 'd1020;
    mem[164] = 'd1020;
    mem[165] = 'd1020;
    mem[166] = 'd1020;
    mem[167] = 'd1020;
    mem[168] = 'd1020;
    mem[169] = 'd1020;
    mem[170] = 'd1020;
    mem[171] = 'd1020;
    mem[172] = 'd1020;
    mem[173] = 'd1020;
    mem[174] = 'd1020;
    mem[175] = 'd1020;
    mem[176] = 'd1020;
    mem[177] = 'd1020;
    mem[178] = 'd1020;
    mem[179] = 'd1020;
    mem[180] = 'd1020;
    mem[181] = 'd1020;
    mem[182] = 'd988;
    mem[183] = 'd1000;
    mem[184] = 'd704;
    mem[185] = 'd872;
    mem[186] = 'd492;
    mem[187] = 'd804;
    mem[188] = 'd340;
    mem[189] = 'd768;
    mem[190] = 'd240;
    mem[191] = 'd748;
    mem[192] = 'd196;
    mem[193] = 'd740;
    mem[194] = 'd196;
    mem[195] = 'd740;
    mem[196] = 'd236;
    mem[197] = 'd744;
    mem[198] = 'd336;
    mem[199] = 'd764;
    mem[200] = 'd480;
    mem[201] = 'd800;
    mem[202] = 'd692;
    mem[203] = 'd868;
    mem[204] = 'd940;
    mem[205] = 'd976;
    mem[206] = 'd1020;
    mem[207] = 'd1020;
    mem[208] = 'd1020;
    mem[209] = 'd1020;
    mem[210] = 'd1020;
    mem[211] = 'd1020;
    mem[212] = 'd1020;
    mem[213] = 'd1020;
    mem[214] = 'd1020;
    mem[215] = 'd1020;
    mem[216] = 'd1020;
    mem[217] = 'd1020;
    mem[218] = 'd1020;
    mem[219] = 'd1020;
    mem[220] = 'd1020;
    mem[221] = 'd1020;
    mem[222] = 'd1020;
    mem[223] = 'd1020;
    mem[224] = 'd1020;
    mem[225] = 'd1020;
    mem[226] = 'd1020;
    mem[227] = 'd1020;
    mem[228] = 'd1020;
    mem[229] = 'd1020;
    mem[230] = 'd1020;
    mem[231] = 'd1020;
    mem[232] = 'd1020;
    mem[233] = 'd1020;
    mem[234] = 'd1020;
    mem[235] = 'd1020;
    mem[236] = 'd1020;
    mem[237] = 'd1020;
    mem[238] = 'd1020;
    mem[239] = 'd1020;
    mem[240] = 'd1020;
    mem[241] = 'd1020;
    mem[242] = 'd1020;
    mem[243] = 'd1020;
    mem[244] = 'd1020;
    mem[245] = 'd1020;
    mem[246] = 'd1020;
    mem[247] = 'd1020;
    mem[248] = 'd1020;
    mem[249] = 'd1020;
    mem[250] = 'd1020;
    mem[251] = 'd1020;
    mem[252] = 'd1020;
    mem[253] = 'd1020;
    mem[254] = 'd1020;
    mem[255] = 'd1020;
    mem[256] = 'd1020;
    mem[257] = 'd1020;
    mem[258] = 'd1020;
    mem[259] = 'd1020;
    mem[260] = 'd1000;
    mem[261] = 'd1012;
    mem[262] = 'd872;
    mem[263] = 'd1000;
    mem[264] = 'd804;
    mem[265] = 'd1000;
    mem[266] = 'd768;
    mem[267] = 'd1000;
    mem[268] = 'd748;
    mem[269] = 'd1000;
    mem[270] = 'd740;
    mem[271] = 'd1000;
    mem[272] = 'd740;
    mem[273] = 'd1000;
    mem[274] = 'd744;
    mem[275] = 'd1000;
    mem[276] = 'd764;
    mem[277] = 'd1000;
    mem[278] = 'd800;
    mem[279] = 'd1000;
    mem[280] = 'd868;
    mem[281] = 'd996;
    mem[282] = 'd976;
    mem[283] = 'd1004;
    mem[284] = 'd1020;
    mem[285] = 'd1020;
    mem[286] = 'd1020;
    mem[287] = 'd1020;
    mem[288] = 'd1020;
    mem[289] = 'd1020;
    mem[290] = 'd1020;
    mem[291] = 'd1020;
    mem[292] = 'd1020;
    mem[293] = 'd1020;
    mem[294] = 'd1020;
    mem[295] = 'd1020;
    mem[296] = 'd1020;
    mem[297] = 'd1020;
    mem[298] = 'd1020;
    mem[299] = 'd1020;
    mem[300] = 'd1020;
    mem[301] = 'd1020;
    mem[302] = 'd1020;
    mem[303] = 'd1020;
    mem[304] = 'd1020;
    mem[305] = 'd1020;
    mem[306] = 'd1020;
    mem[307] = 'd1020;
    mem[308] = 'd1020;
    mem[309] = 'd1020;
    mem[310] = 'd1020;
    mem[311] = 'd1020;
    mem[312] = 'd1020;
    mem[313] = 'd1020;
    mem[314] = 'd1020;
    mem[315] = 'd1020;
    mem[316] = 'd1020;
    mem[317] = 'd1020;
    mem[318] = 'd1020;
    mem[319] = 'd1020;
    mem[320] = 'd1020;
    mem[321] = 'd1020;
    mem[322] = 'd1020;
    mem[323] = 'd1020;
    mem[324] = 'd1020;
    mem[325] = 'd1020;
    mem[326] = 'd1020;
    mem[327] = 'd1020;
    mem[328] = 'd1020;
    mem[329] = 'd1020;
    mem[330] = 'd1020;
    mem[331] = 'd1020;
    mem[332] = 'd1020;
    mem[333] = 'd1020;
    mem[334] = 'd808;
    mem[335] = 'd912;
    mem[336] = 'd408;
    mem[337] = 'd768;
    mem[338] = 'd100;
    mem[339] = 'd696;
    mem[340] = 'd88;
    mem[341] = 'd772;
    mem[342] = 'd96;
    mem[343] = 'd828;
    mem[344] = 'd112;
    mem[345] = 'd868;
    mem[346] = 'd180;
    mem[347] = 'd900;
    mem[348] = 'd224;
    mem[349] = 'd916;
    mem[350] = 'd232;
    mem[351] = 'd916;
    mem[352] = 'd184;
    mem[353] = 'd900;
    mem[354] = 'd120;
    mem[355] = 'd868;
    mem[356] = 'd92;
    mem[357] = 'd828;
    mem[358] = 'd88;
    mem[359] = 'd776;
    mem[360] = 'd128;
    mem[361] = 'd712;
    mem[362] = 'd372;
    mem[363] = 'd752;
    mem[364] = 'd780;
    mem[365] = 'd904;
    mem[366] = 'd1012;
    mem[367] = 'd1012;
    mem[368] = 'd1020;
    mem[369] = 'd1020;
    mem[370] = 'd1020;
    mem[371] = 'd1020;
    mem[372] = 'd1020;
    mem[373] = 'd1020;
    mem[374] = 'd1020;
    mem[375] = 'd1020;
    mem[376] = 'd1020;
    mem[377] = 'd1020;
    mem[378] = 'd1020;
    mem[379] = 'd1020;
    mem[380] = 'd1020;
    mem[381] = 'd1020;
    mem[382] = 'd1020;
    mem[383] = 'd1020;
    mem[384] = 'd1020;
    mem[385] = 'd1020;
    mem[386] = 'd1020;
    mem[387] = 'd1020;
    mem[388] = 'd1020;
    mem[389] = 'd1020;
    mem[390] = 'd1020;
    mem[391] = 'd1020;
    mem[392] = 'd1020;
    mem[393] = 'd1020;
    mem[394] = 'd1020;
    mem[395] = 'd1020;
    mem[396] = 'd1020;
    mem[397] = 'd1020;
    mem[398] = 'd1020;
    mem[399] = 'd1020;
    mem[400] = 'd1020;
    mem[401] = 'd1020;
    mem[402] = 'd1020;
    mem[403] = 'd1020;
    mem[404] = 'd1020;
    mem[405] = 'd1020;
    mem[406] = 'd1020;
    mem[407] = 'd1020;
    mem[408] = 'd1020;
    mem[409] = 'd1020;
    mem[410] = 'd1020;
    mem[411] = 'd1020;
    mem[412] = 'd912;
    mem[413] = 'd996;
    mem[414] = 'd768;
    mem[415] = 'd996;
    mem[416] = 'd696;
    mem[417] = 'd1012;
    mem[418] = 'd772;
    mem[419] = 'd1020;
    mem[420] = 'd828;
    mem[421] = 'd1020;
    mem[422] = 'd868;
    mem[423] = 'd1020;
    mem[424] = 'd900;
    mem[425] = 'd1020;
    mem[426] = 'd916;
    mem[427] = 'd1020;
    mem[428] = 'd916;
    mem[429] = 'd1020;
    mem[430] = 'd900;
    mem[431] = 'd1020;
    mem[432] = 'd868;
    mem[433] = 'd1020;
    mem[434] = 'd828;
    mem[435] = 'd1020;
    mem[436] = 'd776;
    mem[437] = 'd1020;
    mem[438] = 'd712;
    mem[439] = 'd1008;
    mem[440] = 'd752;
    mem[441] = 'd996;
    mem[442] = 'd904;
    mem[443] = 'd1000;
    mem[444] = 'd1012;
    mem[445] = 'd1016;
    mem[446] = 'd1020;
    mem[447] = 'd1020;
    mem[448] = 'd1020;
    mem[449] = 'd1020;
    mem[450] = 'd1020;
    mem[451] = 'd1020;
    mem[452] = 'd1020;
    mem[453] = 'd1020;
    mem[454] = 'd1020;
    mem[455] = 'd1020;
    mem[456] = 'd1020;
    mem[457] = 'd1020;
    mem[458] = 'd1020;
    mem[459] = 'd1020;
    mem[460] = 'd1020;
    mem[461] = 'd1020;
    mem[462] = 'd1020;
    mem[463] = 'd1020;
    mem[464] = 'd1020;
    mem[465] = 'd1020;
    mem[466] = 'd1020;
    mem[467] = 'd1020;
    mem[468] = 'd1020;
    mem[469] = 'd1020;
    mem[470] = 'd1020;
    mem[471] = 'd1020;
    mem[472] = 'd1020;
    mem[473] = 'd1020;
    mem[474] = 'd1020;
    mem[475] = 'd1020;
    mem[476] = 'd1020;
    mem[477] = 'd1020;
    mem[478] = 'd1020;
    mem[479] = 'd1020;
    mem[480] = 'd1020;
    mem[481] = 'd1020;
    mem[482] = 'd1020;
    mem[483] = 'd1020;
    mem[484] = 'd1020;
    mem[485] = 'd1020;
    mem[486] = 'd868;
    mem[487] = 'd936;
    mem[488] = 'd316;
    mem[489] = 'd724;
    mem[490] = 'd52;
    mem[491] = 'd704;
    mem[492] = 'd68;
    mem[493] = 'd792;
    mem[494] = 'd164;
    mem[495] = 'd872;
    mem[496] = 'd480;
    mem[497] = 'd952;
    mem[498] = 'd704;
    mem[499] = 'd992;
    mem[500] = 'd868;
    mem[501] = 'd1012;
    mem[502] = 'd924;
    mem[503] = 'd1016;
    mem[504] = 'd940;
    mem[505] = 'd1016;
    mem[506] = 'd940;
    mem[507] = 'd1016;
    mem[508] = 'd928;
    mem[509] = 'd1016;
    mem[510] = 'd876;
    mem[511] = 'd1012;
    mem[512] = 'd736;
    mem[513] = 'd992;
    mem[514] = 'd516;
    mem[515] = 'd956;
    mem[516] = 'd228;
    mem[517] = 'd876;
    mem[518] = 'd72;
    mem[519] = 'd792;
    mem[520] = 'd64;
    mem[521] = 'd708;
    mem[522] = 'd308;
    mem[523] = 'd724;
    mem[524] = 'd824;
    mem[525] = 'd924;
    mem[526] = 'd1020;
    mem[527] = 'd1020;
    mem[528] = 'd1020;
    mem[529] = 'd1020;
    mem[530] = 'd1020;
    mem[531] = 'd1020;
    mem[532] = 'd1020;
    mem[533] = 'd1020;
    mem[534] = 'd1020;
    mem[535] = 'd1020;
    mem[536] = 'd1020;
    mem[537] = 'd1020;
    mem[538] = 'd1020;
    mem[539] = 'd1020;
    mem[540] = 'd1020;
    mem[541] = 'd1020;
    mem[542] = 'd1020;
    mem[543] = 'd1020;
    mem[544] = 'd1020;
    mem[545] = 'd1020;
    mem[546] = 'd1020;
    mem[547] = 'd1020;
    mem[548] = 'd1020;
    mem[549] = 'd1020;
    mem[550] = 'd1020;
    mem[551] = 'd1020;
    mem[552] = 'd1020;
    mem[553] = 'd1020;
    mem[554] = 'd1020;
    mem[555] = 'd1020;
    mem[556] = 'd1020;
    mem[557] = 'd1020;
    mem[558] = 'd1020;
    mem[559] = 'd1020;
    mem[560] = 'd1020;
    mem[561] = 'd1020;
    mem[562] = 'd1020;
    mem[563] = 'd1020;
    mem[564] = 'd936;
    mem[565] = 'd996;
    mem[566] = 'd724;
    mem[567] = 'd996;
    mem[568] = 'd704;
    mem[569] = 'd1020;
    mem[570] = 'd792;
    mem[571] = 'd1020;
    mem[572] = 'd872;
    mem[573] = 'd1020;
    mem[574] = 'd952;
    mem[575] = 'd1020;
    mem[576] = 'd992;
    mem[577] = 'd1020;
    mem[578] = 'd1012;
    mem[579] = 'd1020;
    mem[580] = 'd1016;
    mem[581] = 'd1020;
    mem[582] = 'd1016;
    mem[583] = 'd1020;
    mem[584] = 'd1016;
    mem[585] = 'd1020;
    mem[586] = 'd1016;
    mem[587] = 'd1020;
    mem[588] = 'd1012;
    mem[589] = 'd1020;
    mem[590] = 'd992;
    mem[591] = 'd1020;
    mem[592] = 'd956;
    mem[593] = 'd1020;
    mem[594] = 'd876;
    mem[595] = 'd1020;
    mem[596] = 'd792;
    mem[597] = 'd1020;
    mem[598] = 'd708;
    mem[599] = 'd1016;
    mem[600] = 'd724;
    mem[601] = 'd996;
    mem[602] = 'd924;
    mem[603] = 'd1000;
    mem[604] = 'd1020;
    mem[605] = 'd1020;
    mem[606] = 'd1020;
    mem[607] = 'd1020;
    mem[608] = 'd1020;
    mem[609] = 'd1020;
    mem[610] = 'd1020;
    mem[611] = 'd1020;
    mem[612] = 'd1020;
    mem[613] = 'd1020;
    mem[614] = 'd1020;
    mem[615] = 'd1020;
    mem[616] = 'd1020;
    mem[617] = 'd1020;
    mem[618] = 'd1020;
    mem[619] = 'd1020;
    mem[620] = 'd1020;
    mem[621] = 'd1020;
    mem[622] = 'd1020;
    mem[623] = 'd1020;
    mem[624] = 'd1020;
    mem[625] = 'd1020;
    mem[626] = 'd1020;
    mem[627] = 'd1020;
    mem[628] = 'd1020;
    mem[629] = 'd1020;
    mem[630] = 'd1020;
    mem[631] = 'd1020;
    mem[632] = 'd1020;
    mem[633] = 'd1020;
    mem[634] = 'd1020;
    mem[635] = 'd1020;
    mem[636] = 'd1020;
    mem[637] = 'd1020;
    mem[638] = 'd1020;
    mem[639] = 'd1020;
    mem[640] = 'd572;
    mem[641] = 'd804;
    mem[642] = 'd52;
    mem[643] = 'd660;
    mem[644] = 'd52;
    mem[645] = 'd764;
    mem[646] = 'd212;
    mem[647] = 'd868;
    mem[648] = 'd600;
    mem[649] = 'd972;
    mem[650] = 'd840;
    mem[651] = 'd1008;
    mem[652] = 'd852;
    mem[653] = 'd1012;
    mem[654] = 'd864;
    mem[655] = 'd1012;
    mem[656] = 'd880;
    mem[657] = 'd1012;
    mem[658] = 'd888;
    mem[659] = 'd1012;
    mem[660] = 'd892;
    mem[661] = 'd1012;
    mem[662] = 'd892;
    mem[663] = 'd1012;
    mem[664] = 'd888;
    mem[665] = 'd1012;
    mem[666] = 'd876;
    mem[667] = 'd1012;
    mem[668] = 'd864;
    mem[669] = 'd1012;
    mem[670] = 'd848;
    mem[671] = 'd1012;
    mem[672] = 'd836;
    mem[673] = 'd1012;
    mem[674] = 'd648;
    mem[675] = 'd976;
    mem[676] = 'd276;
    mem[677] = 'd880;
    mem[678] = 'd60;
    mem[679] = 'd768;
    mem[680] = 'd84;
    mem[681] = 'd680;
    mem[682] = 'd532;
    mem[683] = 'd792;
    mem[684] = 'd988;
    mem[685] = 'd1004;
    mem[686] = 'd1020;
    mem[687] = 'd1020;
    mem[688] = 'd1020;
    mem[689] = 'd1020;
    mem[690] = 'd1020;
    mem[691] = 'd1020;
    mem[692] = 'd1020;
    mem[693] = 'd1020;
    mem[694] = 'd1020;
    mem[695] = 'd1020;
    mem[696] = 'd1020;
    mem[697] = 'd1020;
    mem[698] = 'd1020;
    mem[699] = 'd1020;
    mem[700] = 'd1020;
    mem[701] = 'd1020;
    mem[702] = 'd1020;
    mem[703] = 'd1020;
    mem[704] = 'd1020;
    mem[705] = 'd1020;
    mem[706] = 'd1020;
    mem[707] = 'd1020;
    mem[708] = 'd1020;
    mem[709] = 'd1020;
    mem[710] = 'd1020;
    mem[711] = 'd1020;
    mem[712] = 'd1020;
    mem[713] = 'd1020;
    mem[714] = 'd1020;
    mem[715] = 'd1020;
    mem[716] = 'd1020;
    mem[717] = 'd1020;
    mem[718] = 'd804;
    mem[719] = 'd984;
    mem[720] = 'd660;
    mem[721] = 'd1012;
    mem[722] = 'd764;
    mem[723] = 'd1020;
    mem[724] = 'd868;
    mem[725] = 'd1020;
    mem[726] = 'd972;
    mem[727] = 'd1020;
    mem[728] = 'd1008;
    mem[729] = 'd1020;
    mem[730] = 'd1012;
    mem[731] = 'd1020;
    mem[732] = 'd1012;
    mem[733] = 'd1020;
    mem[734] = 'd1012;
    mem[735] = 'd1020;
    mem[736] = 'd1012;
    mem[737] = 'd1020;
    mem[738] = 'd1012;
    mem[739] = 'd1020;
    mem[740] = 'd1012;
    mem[741] = 'd1020;
    mem[742] = 'd1012;
    mem[743] = 'd1020;
    mem[744] = 'd1012;
    mem[745] = 'd1020;
    mem[746] = 'd1012;
    mem[747] = 'd1020;
    mem[748] = 'd1012;
    mem[749] = 'd1020;
    mem[750] = 'd1012;
    mem[751] = 'd1020;
    mem[752] = 'd976;
    mem[753] = 'd1020;
    mem[754] = 'd880;
    mem[755] = 'd1020;
    mem[756] = 'd768;
    mem[757] = 'd1020;
    mem[758] = 'd680;
    mem[759] = 'd1012;
    mem[760] = 'd792;
    mem[761] = 'd996;
    mem[762] = 'd1004;
    mem[763] = 'd1012;
    mem[764] = 'd1020;
    mem[765] = 'd1020;
    mem[766] = 'd1020;
    mem[767] = 'd1020;
    mem[768] = 'd1020;
    mem[769] = 'd1020;
    mem[770] = 'd1020;
    mem[771] = 'd1020;
    mem[772] = 'd1020;
    mem[773] = 'd1020;
    mem[774] = 'd1020;
    mem[775] = 'd1020;
    mem[776] = 'd1020;
    mem[777] = 'd1020;
    mem[778] = 'd1020;
    mem[779] = 'd1020;
    mem[780] = 'd1020;
    mem[781] = 'd1020;
    mem[782] = 'd1020;
    mem[783] = 'd1020;
    mem[784] = 'd1020;
    mem[785] = 'd1020;
    mem[786] = 'd1020;
    mem[787] = 'd1020;
    mem[788] = 'd1020;
    mem[789] = 'd1020;
    mem[790] = 'd1020;
    mem[791] = 'd1020;
    mem[792] = 'd912;
    mem[793] = 'd964;
    mem[794] = 'd296;
    mem[795] = 'd700;
    mem[796] = 'd36;
    mem[797] = 'd696;
    mem[798] = 'd140;
    mem[799] = 'd816;
    mem[800] = 'd520;
    mem[801] = 'd948;
    mem[802] = 'd764;
    mem[803] = 'd1004;
    mem[804] = 'd776;
    mem[805] = 'd1004;
    mem[806] = 'd788;
    mem[807] = 'd1008;
    mem[808] = 'd804;
    mem[809] = 'd1008;
    mem[810] = 'd820;
    mem[811] = 'd1008;
    mem[812] = 'd836;
    mem[813] = 'd1008;
    mem[814] = 'd844;
    mem[815] = 'd1012;
    mem[816] = 'd848;
    mem[817] = 'd1012;
    mem[818] = 'd848;
    mem[819] = 'd1012;
    mem[820] = 'd840;
    mem[821] = 'd1012;
    mem[822] = 'd832;
    mem[823] = 'd1008;
    mem[824] = 'd816;
    mem[825] = 'd1008;
    mem[826] = 'd800;
    mem[827] = 'd1008;
    mem[828] = 'd784;
    mem[829] = 'd1008;
    mem[830] = 'd772;
    mem[831] = 'd1004;
    mem[832] = 'd760;
    mem[833] = 'd1008;
    mem[834] = 'd588;
    mem[835] = 'd964;
    mem[836] = 'd184;
    mem[837] = 'd828;
    mem[838] = 'd36;
    mem[839] = 'd700;
    mem[840] = 'd268;
    mem[841] = 'd688;
    mem[842] = 'd904;
    mem[843] = 'd960;
    mem[844] = 'd1020;
    mem[845] = 'd1020;
    mem[846] = 'd1020;
    mem[847] = 'd1020;
    mem[848] = 'd1020;
    mem[849] = 'd1020;
    mem[850] = 'd1020;
    mem[851] = 'd1020;
    mem[852] = 'd1020;
    mem[853] = 'd1020;
    mem[854] = 'd1020;
    mem[855] = 'd1020;
    mem[856] = 'd1020;
    mem[857] = 'd1020;
    mem[858] = 'd1020;
    mem[859] = 'd1020;
    mem[860] = 'd1020;
    mem[861] = 'd1020;
    mem[862] = 'd1020;
    mem[863] = 'd1020;
    mem[864] = 'd1020;
    mem[865] = 'd1020;
    mem[866] = 'd1020;
    mem[867] = 'd1020;
    mem[868] = 'd1020;
    mem[869] = 'd1020;
    mem[870] = 'd964;
    mem[871] = 'd1012;
    mem[872] = 'd700;
    mem[873] = 'd988;
    mem[874] = 'd696;
    mem[875] = 'd1020;
    mem[876] = 'd816;
    mem[877] = 'd1020;
    mem[878] = 'd948;
    mem[879] = 'd1020;
    mem[880] = 'd1004;
    mem[881] = 'd1020;
    mem[882] = 'd1004;
    mem[883] = 'd1020;
    mem[884] = 'd1008;
    mem[885] = 'd1020;
    mem[886] = 'd1008;
    mem[887] = 'd1020;
    mem[888] = 'd1008;
    mem[889] = 'd1020;
    mem[890] = 'd1008;
    mem[891] = 'd1020;
    mem[892] = 'd1012;
    mem[893] = 'd1020;
    mem[894] = 'd1012;
    mem[895] = 'd1020;
    mem[896] = 'd1012;
    mem[897] = 'd1020;
    mem[898] = 'd1012;
    mem[899] = 'd1020;
    mem[900] = 'd1008;
    mem[901] = 'd1020;
    mem[902] = 'd1008;
    mem[903] = 'd1020;
    mem[904] = 'd1008;
    mem[905] = 'd1020;
    mem[906] = 'd1008;
    mem[907] = 'd1020;
    mem[908] = 'd1004;
    mem[909] = 'd1020;
    mem[910] = 'd1008;
    mem[911] = 'd1020;
    mem[912] = 'd964;
    mem[913] = 'd1020;
    mem[914] = 'd828;
    mem[915] = 'd1020;
    mem[916] = 'd700;
    mem[917] = 'd1020;
    mem[918] = 'd688;
    mem[919] = 'd988;
    mem[920] = 'd960;
    mem[921] = 'd1012;
    mem[922] = 'd1020;
    mem[923] = 'd1020;
    mem[924] = 'd1020;
    mem[925] = 'd1020;
    mem[926] = 'd1020;
    mem[927] = 'd1020;
    mem[928] = 'd1020;
    mem[929] = 'd1020;
    mem[930] = 'd1020;
    mem[931] = 'd1020;
    mem[932] = 'd1020;
    mem[933] = 'd1020;
    mem[934] = 'd1020;
    mem[935] = 'd1020;
    mem[936] = 'd1020;
    mem[937] = 'd1020;
    mem[938] = 'd1020;
    mem[939] = 'd1020;
    mem[940] = 'd1020;
    mem[941] = 'd1020;
    mem[942] = 'd1020;
    mem[943] = 'd1020;
    mem[944] = 'd1020;
    mem[945] = 'd1020;
    mem[946] = 'd912;
    mem[947] = 'd964;
    mem[948] = 'd188;
    mem[949] = 'd648;
    mem[950] = 'd32;
    mem[951] = 'd708;
    mem[952] = 'd220;
    mem[953] = 'd836;
    mem[954] = 'd632;
    mem[955] = 'd976;
    mem[956] = 'd696;
    mem[957] = 'd1004;
    mem[958] = 'd708;
    mem[959] = 'd1004;
    mem[960] = 'd720;
    mem[961] = 'd1004;
    mem[962] = 'd736;
    mem[963] = 'd1004;
    mem[964] = 'd752;
    mem[965] = 'd1004;
    mem[966] = 'd764;
    mem[967] = 'd1004;
    mem[968] = 'd780;
    mem[969] = 'd1004;
    mem[970] = 'd788;
    mem[971] = 'd1008;
    mem[972] = 'd796;
    mem[973] = 'd1008;
    mem[974] = 'd792;
    mem[975] = 'd1008;
    mem[976] = 'd788;
    mem[977] = 'd1004;
    mem[978] = 'd780;
    mem[979] = 'd1004;
    mem[980] = 'd764;
    mem[981] = 'd1004;
    mem[982] = 'd748;
    mem[983] = 'd1004;
    mem[984] = 'd732;
    mem[985] = 'd1004;
    mem[986] = 'd716;
    mem[987] = 'd1004;
    mem[988] = 'd704;
    mem[989] = 'd1004;
    mem[990] = 'd692;
    mem[991] = 'd1004;
    mem[992] = 'd656;
    mem[993] = 'd980;
    mem[994] = 'd300;
    mem[995] = 'd860;
    mem[996] = 'd32;
    mem[997] = 'd708;
    mem[998] = 'd160;
    mem[999] = 'd644;
    mem[1000] = 'd904;
    mem[1001] = 'd960;
    mem[1002] = 'd1020;
    mem[1003] = 'd1020;
    mem[1004] = 'd1020;
    mem[1005] = 'd1020;
    mem[1006] = 'd1020;
    mem[1007] = 'd1020;
    mem[1008] = 'd1020;
    mem[1009] = 'd1020;
    mem[1010] = 'd1020;
    mem[1011] = 'd1020;
    mem[1012] = 'd1020;
    mem[1013] = 'd1020;
    mem[1014] = 'd1020;
    mem[1015] = 'd1020;
    mem[1016] = 'd1020;
    mem[1017] = 'd1020;
    mem[1018] = 'd1020;
    mem[1019] = 'd1020;
    mem[1020] = 'd1020;
    mem[1021] = 'd1020;
    mem[1022] = 'd1020;
    mem[1023] = 'd1020;
    mem[1024] = 'd964;
    mem[1025] = 'd1008;
    mem[1026] = 'd648;
    mem[1027] = 'd992;
    mem[1028] = 'd708;
    mem[1029] = 'd1020;
    mem[1030] = 'd836;
    mem[1031] = 'd1020;
    mem[1032] = 'd976;
    mem[1033] = 'd1020;
    mem[1034] = 'd1004;
    mem[1035] = 'd1020;
    mem[1036] = 'd1004;
    mem[1037] = 'd1020;
    mem[1038] = 'd1004;
    mem[1039] = 'd1020;
    mem[1040] = 'd1004;
    mem[1041] = 'd1020;
    mem[1042] = 'd1004;
    mem[1043] = 'd1020;
    mem[1044] = 'd1004;
    mem[1045] = 'd1020;
    mem[1046] = 'd1004;
    mem[1047] = 'd1020;
    mem[1048] = 'd1008;
    mem[1049] = 'd1020;
    mem[1050] = 'd1008;
    mem[1051] = 'd1020;
    mem[1052] = 'd1008;
    mem[1053] = 'd1020;
    mem[1054] = 'd1004;
    mem[1055] = 'd1020;
    mem[1056] = 'd1004;
    mem[1057] = 'd1020;
    mem[1058] = 'd1004;
    mem[1059] = 'd1020;
    mem[1060] = 'd1004;
    mem[1061] = 'd1020;
    mem[1062] = 'd1004;
    mem[1063] = 'd1020;
    mem[1064] = 'd1004;
    mem[1065] = 'd1020;
    mem[1066] = 'd1004;
    mem[1067] = 'd1020;
    mem[1068] = 'd1004;
    mem[1069] = 'd1020;
    mem[1070] = 'd980;
    mem[1071] = 'd1020;
    mem[1072] = 'd860;
    mem[1073] = 'd1020;
    mem[1074] = 'd708;
    mem[1075] = 'd1020;
    mem[1076] = 'd644;
    mem[1077] = 'd996;
    mem[1078] = 'd960;
    mem[1079] = 'd1012;
    mem[1080] = 'd1020;
    mem[1081] = 'd1020;
    mem[1082] = 'd1020;
    mem[1083] = 'd1020;
    mem[1084] = 'd1020;
    mem[1085] = 'd1020;
    mem[1086] = 'd1020;
    mem[1087] = 'd1020;
    mem[1088] = 'd1020;
    mem[1089] = 'd1020;
    mem[1090] = 'd1020;
    mem[1091] = 'd1020;
    mem[1092] = 'd1020;
    mem[1093] = 'd1020;
    mem[1094] = 'd1020;
    mem[1095] = 'd1020;
    mem[1096] = 'd1020;
    mem[1097] = 'd1020;
    mem[1098] = 'd1020;
    mem[1099] = 'd1020;
    mem[1100] = 'd964;
    mem[1101] = 'd984;
    mem[1102] = 'd248;
    mem[1103] = 'd660;
    mem[1104] = 'd32;
    mem[1105] = 'd688;
    mem[1106] = 'd232;
    mem[1107] = 'd832;
    mem[1108] = 'd592;
    mem[1109] = 'd960;
    mem[1110] = 'd628;
    mem[1111] = 'd988;
    mem[1112] = 'd640;
    mem[1113] = 'd996;
    mem[1114] = 'd652;
    mem[1115] = 'd1000;
    mem[1116] = 'd664;
    mem[1117] = 'd1000;
    mem[1118] = 'd676;
    mem[1119] = 'd1000;
    mem[1120] = 'd692;
    mem[1121] = 'd1004;
    mem[1122] = 'd708;
    mem[1123] = 'd1004;
    mem[1124] = 'd716;
    mem[1125] = 'd1004;
    mem[1126] = 'd728;
    mem[1127] = 'd1004;
    mem[1128] = 'd732;
    mem[1129] = 'd1004;
    mem[1130] = 'd732;
    mem[1131] = 'd1004;
    mem[1132] = 'd724;
    mem[1133] = 'd1004;
    mem[1134] = 'd716;
    mem[1135] = 'd1004;
    mem[1136] = 'd704;
    mem[1137] = 'd1004;
    mem[1138] = 'd692;
    mem[1139] = 'd1004;
    mem[1140] = 'd676;
    mem[1141] = 'd1000;
    mem[1142] = 'd664;
    mem[1143] = 'd1000;
    mem[1144] = 'd652;
    mem[1145] = 'd1000;
    mem[1146] = 'd640;
    mem[1147] = 'd996;
    mem[1148] = 'd628;
    mem[1149] = 'd988;
    mem[1150] = 'd616;
    mem[1151] = 'd964;
    mem[1152] = 'd300;
    mem[1153] = 'd852;
    mem[1154] = 'd28;
    mem[1155] = 'd692;
    mem[1156] = 'd212;
    mem[1157] = 'd648;
    mem[1158] = 'd948;
    mem[1159] = 'd976;
    mem[1160] = 'd1020;
    mem[1161] = 'd1020;
    mem[1162] = 'd1020;
    mem[1163] = 'd1020;
    mem[1164] = 'd1020;
    mem[1165] = 'd1020;
    mem[1166] = 'd1020;
    mem[1167] = 'd1020;
    mem[1168] = 'd1020;
    mem[1169] = 'd1020;
    mem[1170] = 'd1020;
    mem[1171] = 'd1020;
    mem[1172] = 'd1020;
    mem[1173] = 'd1020;
    mem[1174] = 'd1020;
    mem[1175] = 'd1020;
    mem[1176] = 'd1020;
    mem[1177] = 'd1020;
    mem[1178] = 'd984;
    mem[1179] = 'd1004;
    mem[1180] = 'd660;
    mem[1181] = 'd980;
    mem[1182] = 'd688;
    mem[1183] = 'd1020;
    mem[1184] = 'd832;
    mem[1185] = 'd1020;
    mem[1186] = 'd960;
    mem[1187] = 'd1020;
    mem[1188] = 'd988;
    mem[1189] = 'd1020;
    mem[1190] = 'd996;
    mem[1191] = 'd1020;
    mem[1192] = 'd1000;
    mem[1193] = 'd1020;
    mem[1194] = 'd1000;
    mem[1195] = 'd1020;
    mem[1196] = 'd1000;
    mem[1197] = 'd1020;
    mem[1198] = 'd1004;
    mem[1199] = 'd1020;
    mem[1200] = 'd1004;
    mem[1201] = 'd1020;
    mem[1202] = 'd1004;
    mem[1203] = 'd1020;
    mem[1204] = 'd1004;
    mem[1205] = 'd1020;
    mem[1206] = 'd1004;
    mem[1207] = 'd1020;
    mem[1208] = 'd1004;
    mem[1209] = 'd1020;
    mem[1210] = 'd1004;
    mem[1211] = 'd1020;
    mem[1212] = 'd1004;
    mem[1213] = 'd1020;
    mem[1214] = 'd1004;
    mem[1215] = 'd1020;
    mem[1216] = 'd1004;
    mem[1217] = 'd1020;
    mem[1218] = 'd1000;
    mem[1219] = 'd1020;
    mem[1220] = 'd1000;
    mem[1221] = 'd1020;
    mem[1222] = 'd1000;
    mem[1223] = 'd1020;
    mem[1224] = 'd996;
    mem[1225] = 'd1020;
    mem[1226] = 'd988;
    mem[1227] = 'd1020;
    mem[1228] = 'd964;
    mem[1229] = 'd1020;
    mem[1230] = 'd852;
    mem[1231] = 'd1020;
    mem[1232] = 'd692;
    mem[1233] = 'd1020;
    mem[1234] = 'd648;
    mem[1235] = 'd984;
    mem[1236] = 'd976;
    mem[1237] = 'd1004;
    mem[1238] = 'd1020;
    mem[1239] = 'd1020;
    mem[1240] = 'd1020;
    mem[1241] = 'd1020;
    mem[1242] = 'd1020;
    mem[1243] = 'd1020;
    mem[1244] = 'd1020;
    mem[1245] = 'd1020;
    mem[1246] = 'd1020;
    mem[1247] = 'd1020;
    mem[1248] = 'd1020;
    mem[1249] = 'd1020;
    mem[1250] = 'd1020;
    mem[1251] = 'd1020;
    mem[1252] = 'd1020;
    mem[1253] = 'd1020;
    mem[1254] = 'd1020;
    mem[1255] = 'd1020;
    mem[1256] = 'd452;
    mem[1257] = 'd748;
    mem[1258] = 'd24;
    mem[1259] = 'd656;
    mem[1260] = 'd160;
    mem[1261] = 'd796;
    mem[1262] = 'd524;
    mem[1263] = 'd932;
    mem[1264] = 'd560;
    mem[1265] = 'd964;
    mem[1266] = 'd572;
    mem[1267] = 'd984;
    mem[1268] = 'd584;
    mem[1269] = 'd996;
    mem[1270] = 'd592;
    mem[1271] = 'd996;
    mem[1272] = 'd604;
    mem[1273] = 'd996;
    mem[1274] = 'd616;
    mem[1275] = 'd996;
    mem[1276] = 'd628;
    mem[1277] = 'd996;
    mem[1278] = 'd644;
    mem[1279] = 'd1000;
    mem[1280] = 'd652;
    mem[1281] = 'd1000;
    mem[1282] = 'd660;
    mem[1283] = 'd1000;
    mem[1284] = 'd664;
    mem[1285] = 'd1000;
    mem[1286] = 'd664;
    mem[1287] = 'd1000;
    mem[1288] = 'd660;
    mem[1289] = 'd1000;
    mem[1290] = 'd652;
    mem[1291] = 'd1000;
    mem[1292] = 'd640;
    mem[1293] = 'd1000;
    mem[1294] = 'd628;
    mem[1295] = 'd996;
    mem[1296] = 'd616;
    mem[1297] = 'd996;
    mem[1298] = 'd604;
    mem[1299] = 'd996;
    mem[1300] = 'd592;
    mem[1301] = 'd996;
    mem[1302] = 'd584;
    mem[1303] = 'd996;
    mem[1304] = 'd572;
    mem[1305] = 'd988;
    mem[1306] = 'd560;
    mem[1307] = 'd968;
    mem[1308] = 'd544;
    mem[1309] = 'd936;
    mem[1310] = 'd232;
    mem[1311] = 'd812;
    mem[1312] = 'd24;
    mem[1313] = 'd660;
    mem[1314] = 'd468;
    mem[1315] = 'd752;
    mem[1316] = 'd1020;
    mem[1317] = 'd1020;
    mem[1318] = 'd1020;
    mem[1319] = 'd1020;
    mem[1320] = 'd1020;
    mem[1321] = 'd1020;
    mem[1322] = 'd1020;
    mem[1323] = 'd1020;
    mem[1324] = 'd1020;
    mem[1325] = 'd1020;
    mem[1326] = 'd1020;
    mem[1327] = 'd1020;
    mem[1328] = 'd1020;
    mem[1329] = 'd1020;
    mem[1330] = 'd1020;
    mem[1331] = 'd1020;
    mem[1332] = 'd1020;
    mem[1333] = 'd1020;
    mem[1334] = 'd748;
    mem[1335] = 'd988;
    mem[1336] = 'd656;
    mem[1337] = 'd1020;
    mem[1338] = 'd796;
    mem[1339] = 'd1020;
    mem[1340] = 'd932;
    mem[1341] = 'd1020;
    mem[1342] = 'd964;
    mem[1343] = 'd1020;
    mem[1344] = 'd984;
    mem[1345] = 'd1020;
    mem[1346] = 'd996;
    mem[1347] = 'd1020;
    mem[1348] = 'd996;
    mem[1349] = 'd1020;
    mem[1350] = 'd996;
    mem[1351] = 'd1020;
    mem[1352] = 'd996;
    mem[1353] = 'd1020;
    mem[1354] = 'd996;
    mem[1355] = 'd1020;
    mem[1356] = 'd1000;
    mem[1357] = 'd1020;
    mem[1358] = 'd1000;
    mem[1359] = 'd1020;
    mem[1360] = 'd1000;
    mem[1361] = 'd1020;
    mem[1362] = 'd1000;
    mem[1363] = 'd1020;
    mem[1364] = 'd1000;
    mem[1365] = 'd1020;
    mem[1366] = 'd1000;
    mem[1367] = 'd1020;
    mem[1368] = 'd1000;
    mem[1369] = 'd1020;
    mem[1370] = 'd1000;
    mem[1371] = 'd1020;
    mem[1372] = 'd996;
    mem[1373] = 'd1020;
    mem[1374] = 'd996;
    mem[1375] = 'd1020;
    mem[1376] = 'd996;
    mem[1377] = 'd1020;
    mem[1378] = 'd996;
    mem[1379] = 'd1020;
    mem[1380] = 'd996;
    mem[1381] = 'd1020;
    mem[1382] = 'd988;
    mem[1383] = 'd1020;
    mem[1384] = 'd968;
    mem[1385] = 'd1020;
    mem[1386] = 'd936;
    mem[1387] = 'd1020;
    mem[1388] = 'd812;
    mem[1389] = 'd1020;
    mem[1390] = 'd660;
    mem[1391] = 'd1020;
    mem[1392] = 'd752;
    mem[1393] = 'd984;
    mem[1394] = 'd1020;
    mem[1395] = 'd1020;
    mem[1396] = 'd1020;
    mem[1397] = 'd1020;
    mem[1398] = 'd1020;
    mem[1399] = 'd1020;
    mem[1400] = 'd1020;
    mem[1401] = 'd1020;
    mem[1402] = 'd1020;
    mem[1403] = 'd1020;
    mem[1404] = 'd1020;
    mem[1405] = 'd1020;
    mem[1406] = 'd1020;
    mem[1407] = 'd1020;
    mem[1408] = 'd1020;
    mem[1409] = 'd1020;
    mem[1410] = 'd840;
    mem[1411] = 'd924;
    mem[1412] = 'd32;
    mem[1413] = 'd608;
    mem[1414] = 'd76;
    mem[1415] = 'd736;
    mem[1416] = 'd436;
    mem[1417] = 'd896;
    mem[1418] = 'd496;
    mem[1419] = 'd936;
    mem[1420] = 'd508;
    mem[1421] = 'd956;
    mem[1422] = 'd516;
    mem[1423] = 'd976;
    mem[1424] = 'd528;
    mem[1425] = 'd992;
    mem[1426] = 'd536;
    mem[1427] = 'd992;
    mem[1428] = 'd544;
    mem[1429] = 'd996;
    mem[1430] = 'd556;
    mem[1431] = 'd996;
    mem[1432] = 'd568;
    mem[1433] = 'd996;
    mem[1434] = 'd576;
    mem[1435] = 'd996;
    mem[1436] = 'd584;
    mem[1437] = 'd996;
    mem[1438] = 'd592;
    mem[1439] = 'd996;
    mem[1440] = 'd596;
    mem[1441] = 'd996;
    mem[1442] = 'd596;
    mem[1443] = 'd996;
    mem[1444] = 'd592;
    mem[1445] = 'd996;
    mem[1446] = 'd584;
    mem[1447] = 'd996;
    mem[1448] = 'd576;
    mem[1449] = 'd996;
    mem[1450] = 'd564;
    mem[1451] = 'd996;
    mem[1452] = 'd556;
    mem[1453] = 'd996;
    mem[1454] = 'd544;
    mem[1455] = 'd996;
    mem[1456] = 'd532;
    mem[1457] = 'd992;
    mem[1458] = 'd524;
    mem[1459] = 'd992;
    mem[1460] = 'd516;
    mem[1461] = 'd976;
    mem[1462] = 'd508;
    mem[1463] = 'd956;
    mem[1464] = 'd496;
    mem[1465] = 'd936;
    mem[1466] = 'd460;
    mem[1467] = 'd900;
    mem[1468] = 'd116;
    mem[1469] = 'd748;
    mem[1470] = 'd28;
    mem[1471] = 'd604;
    mem[1472] = 'd828;
    mem[1473] = 'd912;
    mem[1474] = 'd1020;
    mem[1475] = 'd1020;
    mem[1476] = 'd1020;
    mem[1477] = 'd1020;
    mem[1478] = 'd1020;
    mem[1479] = 'd1020;
    mem[1480] = 'd1020;
    mem[1481] = 'd1020;
    mem[1482] = 'd1020;
    mem[1483] = 'd1020;
    mem[1484] = 'd1020;
    mem[1485] = 'd1020;
    mem[1486] = 'd1020;
    mem[1487] = 'd1020;
    mem[1488] = 'd924;
    mem[1489] = 'd996;
    mem[1490] = 'd608;
    mem[1491] = 'd1008;
    mem[1492] = 'd736;
    mem[1493] = 'd1020;
    mem[1494] = 'd896;
    mem[1495] = 'd1020;
    mem[1496] = 'd936;
    mem[1497] = 'd1020;
    mem[1498] = 'd956;
    mem[1499] = 'd1020;
    mem[1500] = 'd976;
    mem[1501] = 'd1020;
    mem[1502] = 'd992;
    mem[1503] = 'd1020;
    mem[1504] = 'd992;
    mem[1505] = 'd1020;
    mem[1506] = 'd996;
    mem[1507] = 'd1020;
    mem[1508] = 'd996;
    mem[1509] = 'd1020;
    mem[1510] = 'd996;
    mem[1511] = 'd1020;
    mem[1512] = 'd996;
    mem[1513] = 'd1020;
    mem[1514] = 'd996;
    mem[1515] = 'd1020;
    mem[1516] = 'd996;
    mem[1517] = 'd1020;
    mem[1518] = 'd996;
    mem[1519] = 'd1020;
    mem[1520] = 'd996;
    mem[1521] = 'd1020;
    mem[1522] = 'd996;
    mem[1523] = 'd1020;
    mem[1524] = 'd996;
    mem[1525] = 'd1020;
    mem[1526] = 'd996;
    mem[1527] = 'd1020;
    mem[1528] = 'd996;
    mem[1529] = 'd1020;
    mem[1530] = 'd996;
    mem[1531] = 'd1020;
    mem[1532] = 'd996;
    mem[1533] = 'd1020;
    mem[1534] = 'd992;
    mem[1535] = 'd1020;
    mem[1536] = 'd992;
    mem[1537] = 'd1020;
    mem[1538] = 'd976;
    mem[1539] = 'd1020;
    mem[1540] = 'd956;
    mem[1541] = 'd1020;
    mem[1542] = 'd936;
    mem[1543] = 'd1020;
    mem[1544] = 'd900;
    mem[1545] = 'd1020;
    mem[1546] = 'd748;
    mem[1547] = 'd1020;
    mem[1548] = 'd604;
    mem[1549] = 'd1012;
    mem[1550] = 'd912;
    mem[1551] = 'd988;
    mem[1552] = 'd1020;
    mem[1553] = 'd1020;
    mem[1554] = 'd1020;
    mem[1555] = 'd1020;
    mem[1556] = 'd1020;
    mem[1557] = 'd1020;
    mem[1558] = 'd1020;
    mem[1559] = 'd1020;
    mem[1560] = 'd1020;
    mem[1561] = 'd1020;
    mem[1562] = 'd1020;
    mem[1563] = 'd1020;
    mem[1564] = 'd1012;
    mem[1565] = 'd1016;
    mem[1566] = 'd304;
    mem[1567] = 'd668;
    mem[1568] = 'd32;
    mem[1569] = 'd668;
    mem[1570] = 'd284;
    mem[1571] = 'd824;
    mem[1572] = 'd428;
    mem[1573] = 'd900;
    mem[1574] = 'd440;
    mem[1575] = 'd924;
    mem[1576] = 'd452;
    mem[1577] = 'd948;
    mem[1578] = 'd456;
    mem[1579] = 'd964;
    mem[1580] = 'd464;
    mem[1581] = 'd976;
    mem[1582] = 'd476;
    mem[1583] = 'd988;
    mem[1584] = 'd484;
    mem[1585] = 'd988;
    mem[1586] = 'd492;
    mem[1587] = 'd988;
    mem[1588] = 'd504;
    mem[1589] = 'd992;
    mem[1590] = 'd512;
    mem[1591] = 'd992;
    mem[1592] = 'd520;
    mem[1593] = 'd992;
    mem[1594] = 'd524;
    mem[1595] = 'd992;
    mem[1596] = 'd528;
    mem[1597] = 'd992;
    mem[1598] = 'd528;
    mem[1599] = 'd992;
    mem[1600] = 'd524;
    mem[1601] = 'd992;
    mem[1602] = 'd520;
    mem[1603] = 'd992;
    mem[1604] = 'd508;
    mem[1605] = 'd992;
    mem[1606] = 'd504;
    mem[1607] = 'd992;
    mem[1608] = 'd492;
    mem[1609] = 'd988;
    mem[1610] = 'd484;
    mem[1611] = 'd988;
    mem[1612] = 'd476;
    mem[1613] = 'd988;
    mem[1614] = 'd464;
    mem[1615] = 'd976;
    mem[1616] = 'd460;
    mem[1617] = 'd964;
    mem[1618] = 'd448;
    mem[1619] = 'd948;
    mem[1620] = 'd440;
    mem[1621] = 'd928;
    mem[1622] = 'd428;
    mem[1623] = 'd900;
    mem[1624] = 'd336;
    mem[1625] = 'd844;
    mem[1626] = 'd40;
    mem[1627] = 'd672;
    mem[1628] = 'd256;
    mem[1629] = 'd644;
    mem[1630] = 'd1020;
    mem[1631] = 'd1020;
    mem[1632] = 'd1020;
    mem[1633] = 'd1020;
    mem[1634] = 'd1020;
    mem[1635] = 'd1020;
    mem[1636] = 'd1020;
    mem[1637] = 'd1020;
    mem[1638] = 'd1020;
    mem[1639] = 'd1020;
    mem[1640] = 'd1020;
    mem[1641] = 'd1020;
    mem[1642] = 'd1016;
    mem[1643] = 'd1016;
    mem[1644] = 'd668;
    mem[1645] = 'd972;
    mem[1646] = 'd668;
    mem[1647] = 'd1020;
    mem[1648] = 'd824;
    mem[1649] = 'd1020;
    mem[1650] = 'd900;
    mem[1651] = 'd1020;
    mem[1652] = 'd924;
    mem[1653] = 'd1020;
    mem[1654] = 'd948;
    mem[1655] = 'd1020;
    mem[1656] = 'd964;
    mem[1657] = 'd1020;
    mem[1658] = 'd976;
    mem[1659] = 'd1020;
    mem[1660] = 'd988;
    mem[1661] = 'd1020;
    mem[1662] = 'd988;
    mem[1663] = 'd1020;
    mem[1664] = 'd988;
    mem[1665] = 'd1020;
    mem[1666] = 'd992;
    mem[1667] = 'd1020;
    mem[1668] = 'd992;
    mem[1669] = 'd1020;
    mem[1670] = 'd992;
    mem[1671] = 'd1020;
    mem[1672] = 'd992;
    mem[1673] = 'd1020;
    mem[1674] = 'd992;
    mem[1675] = 'd1020;
    mem[1676] = 'd992;
    mem[1677] = 'd1020;
    mem[1678] = 'd992;
    mem[1679] = 'd1020;
    mem[1680] = 'd992;
    mem[1681] = 'd1020;
    mem[1682] = 'd992;
    mem[1683] = 'd1020;
    mem[1684] = 'd992;
    mem[1685] = 'd1020;
    mem[1686] = 'd988;
    mem[1687] = 'd1020;
    mem[1688] = 'd988;
    mem[1689] = 'd1020;
    mem[1690] = 'd988;
    mem[1691] = 'd1020;
    mem[1692] = 'd976;
    mem[1693] = 'd1020;
    mem[1694] = 'd964;
    mem[1695] = 'd1020;
    mem[1696] = 'd948;
    mem[1697] = 'd1020;
    mem[1698] = 'd928;
    mem[1699] = 'd1020;
    mem[1700] = 'd900;
    mem[1701] = 'd1020;
    mem[1702] = 'd844;
    mem[1703] = 'd1020;
    mem[1704] = 'd672;
    mem[1705] = 'd1020;
    mem[1706] = 'd644;
    mem[1707] = 'd972;
    mem[1708] = 'd1020;
    mem[1709] = 'd1020;
    mem[1710] = 'd1020;
    mem[1711] = 'd1020;
    mem[1712] = 'd1020;
    mem[1713] = 'd1020;
    mem[1714] = 'd1020;
    mem[1715] = 'd1020;
    mem[1716] = 'd1020;
    mem[1717] = 'd1020;
    mem[1718] = 'd1020;
    mem[1719] = 'd1020;
    mem[1720] = 'd788;
    mem[1721] = 'd892;
    mem[1722] = 'd24;
    mem[1723] = 'd584;
    mem[1724] = 'd108;
    mem[1725] = 'd700;
    mem[1726] = 'd344;
    mem[1727] = 'd804;
    mem[1728] = 'd356;
    mem[1729] = 'd824;
    mem[1730] = 'd364;
    mem[1731] = 'd840;
    mem[1732] = 'd372;
    mem[1733] = 'd860;
    mem[1734] = 'd388;
    mem[1735] = 'd888;
    mem[1736] = 'd396;
    mem[1737] = 'd912;
    mem[1738] = 'd408;
    mem[1739] = 'd952;
    mem[1740] = 'd424;
    mem[1741] = 'd988;
    mem[1742] = 'd436;
    mem[1743] = 'd992;
    mem[1744] = 'd436;
    mem[1745] = 'd988;
    mem[1746] = 'd448;
    mem[1747] = 'd988;
    mem[1748] = 'd456;
    mem[1749] = 'd988;
    mem[1750] = 'd456;
    mem[1751] = 'd988;
    mem[1752] = 'd460;
    mem[1753] = 'd988;
    mem[1754] = 'd460;
    mem[1755] = 'd988;
    mem[1756] = 'd460;
    mem[1757] = 'd988;
    mem[1758] = 'd456;
    mem[1759] = 'd988;
    mem[1760] = 'd444;
    mem[1761] = 'd988;
    mem[1762] = 'd436;
    mem[1763] = 'd992;
    mem[1764] = 'd432;
    mem[1765] = 'd992;
    mem[1766] = 'd424;
    mem[1767] = 'd980;
    mem[1768] = 'd404;
    mem[1769] = 'd944;
    mem[1770] = 'd392;
    mem[1771] = 'd908;
    mem[1772] = 'd380;
    mem[1773] = 'd884;
    mem[1774] = 'd376;
    mem[1775] = 'd860;
    mem[1776] = 'd368;
    mem[1777] = 'd844;
    mem[1778] = 'd356;
    mem[1779] = 'd828;
    mem[1780] = 'd348;
    mem[1781] = 'd812;
    mem[1782] = 'd148;
    mem[1783] = 'd728;
    mem[1784] = 'd16;
    mem[1785] = 'd584;
    mem[1786] = 'd760;
    mem[1787] = 'd872;
    mem[1788] = 'd1020;
    mem[1789] = 'd1020;
    mem[1790] = 'd1020;
    mem[1791] = 'd1020;
    mem[1792] = 'd1020;
    mem[1793] = 'd1020;
    mem[1794] = 'd1020;
    mem[1795] = 'd1020;
    mem[1796] = 'd1020;
    mem[1797] = 'd1020;
    mem[1798] = 'd892;
    mem[1799] = 'd984;
    mem[1800] = 'd584;
    mem[1801] = 'd1000;
    mem[1802] = 'd700;
    mem[1803] = 'd968;
    mem[1804] = 'd804;
    mem[1805] = 'd948;
    mem[1806] = 'd824;
    mem[1807] = 'd940;
    mem[1808] = 'd840;
    mem[1809] = 'd932;
    mem[1810] = 'd860;
    mem[1811] = 'd936;
    mem[1812] = 'd888;
    mem[1813] = 'd944;
    mem[1814] = 'd912;
    mem[1815] = 'd956;
    mem[1816] = 'd952;
    mem[1817] = 'd980;
    mem[1818] = 'd988;
    mem[1819] = 'd1012;
    mem[1820] = 'd992;
    mem[1821] = 'd1020;
    mem[1822] = 'd988;
    mem[1823] = 'd1020;
    mem[1824] = 'd988;
    mem[1825] = 'd1020;
    mem[1826] = 'd988;
    mem[1827] = 'd1020;
    mem[1828] = 'd988;
    mem[1829] = 'd1020;
    mem[1830] = 'd988;
    mem[1831] = 'd1020;
    mem[1832] = 'd988;
    mem[1833] = 'd1020;
    mem[1834] = 'd988;
    mem[1835] = 'd1020;
    mem[1836] = 'd988;
    mem[1837] = 'd1020;
    mem[1838] = 'd988;
    mem[1839] = 'd1020;
    mem[1840] = 'd992;
    mem[1841] = 'd1020;
    mem[1842] = 'd992;
    mem[1843] = 'd1020;
    mem[1844] = 'd980;
    mem[1845] = 'd1008;
    mem[1846] = 'd944;
    mem[1847] = 'd976;
    mem[1848] = 'd908;
    mem[1849] = 'd956;
    mem[1850] = 'd884;
    mem[1851] = 'd940;
    mem[1852] = 'd860;
    mem[1853] = 'd932;
    mem[1854] = 'd844;
    mem[1855] = 'd936;
    mem[1856] = 'd828;
    mem[1857] = 'd940;
    mem[1858] = 'd812;
    mem[1859] = 'd952;
    mem[1860] = 'd728;
    mem[1861] = 'd988;
    mem[1862] = 'd584;
    mem[1863] = 'd1004;
    mem[1864] = 'd872;
    mem[1865] = 'd976;
    mem[1866] = 'd1020;
    mem[1867] = 'd1020;
    mem[1868] = 'd1020;
    mem[1869] = 'd1020;
    mem[1870] = 'd1020;
    mem[1871] = 'd1020;
    mem[1872] = 'd1020;
    mem[1873] = 'd1020;
    mem[1874] = 'd1020;
    mem[1875] = 'd1020;
    mem[1876] = 'd352;
    mem[1877] = 'd676;
    mem[1878] = 'd52;
    mem[1879] = 'd460;
    mem[1880] = 'd132;
    mem[1881] = 'd168;
    mem[1882] = 'd152;
    mem[1883] = 'd168;
    mem[1884] = 'd152;
    mem[1885] = 'd168;
    mem[1886] = 'd148;
    mem[1887] = 'd160;
    mem[1888] = 'd140;
    mem[1889] = 'd152;
    mem[1890] = 'd144;
    mem[1891] = 'd160;
    mem[1892] = 'd152;
    mem[1893] = 'd176;
    mem[1894] = 'd172;
    mem[1895] = 'd220;
    mem[1896] = 'd204;
    mem[1897] = 'd304;
    mem[1898] = 'd248;
    mem[1899] = 'd428;
    mem[1900] = 'd308;
    mem[1901] = 'd628;
    mem[1902] = 'd340;
    mem[1903] = 'd820;
    mem[1904] = 'd392;
    mem[1905] = 'd980;
    mem[1906] = 'd396;
    mem[1907] = 'd988;
    mem[1908] = 'd396;
    mem[1909] = 'd984;
    mem[1910] = 'd396;
    mem[1911] = 'd988;
    mem[1912] = 'd396;
    mem[1913] = 'd988;
    mem[1914] = 'd380;
    mem[1915] = 'd944;
    mem[1916] = 'd336;
    mem[1917] = 'd788;
    mem[1918] = 'd296;
    mem[1919] = 'd596;
    mem[1920] = 'd244;
    mem[1921] = 'd408;
    mem[1922] = 'd200;
    mem[1923] = 'd288;
    mem[1924] = 'd172;
    mem[1925] = 'd212;
    mem[1926] = 'd152;
    mem[1927] = 'd172;
    mem[1928] = 'd144;
    mem[1929] = 'd164;
    mem[1930] = 'd144;
    mem[1931] = 'd156;
    mem[1932] = 'd156;
    mem[1933] = 'd168;
    mem[1934] = 'd156;
    mem[1935] = 'd172;
    mem[1936] = 'd152;
    mem[1937] = 'd172;
    mem[1938] = 'd132;
    mem[1939] = 'd168;
    mem[1940] = 'd44;
    mem[1941] = 'd540;
    mem[1942] = 'd332;
    mem[1943] = 'd668;
    mem[1944] = 'd1020;
    mem[1945] = 'd1020;
    mem[1946] = 'd1020;
    mem[1947] = 'd1020;
    mem[1948] = 'd1020;
    mem[1949] = 'd1020;
    mem[1950] = 'd1020;
    mem[1951] = 'd1020;
    mem[1952] = 'd1020;
    mem[1953] = 'd1020;
    mem[1954] = 'd676;
    mem[1955] = 'd952;
    mem[1956] = 'd460;
    mem[1957] = 'd732;
    mem[1958] = 'd168;
    mem[1959] = 'd184;
    mem[1960] = 'd168;
    mem[1961] = 'd172;
    mem[1962] = 'd168;
    mem[1963] = 'd168;
    mem[1964] = 'd160;
    mem[1965] = 'd160;
    mem[1966] = 'd152;
    mem[1967] = 'd156;
    mem[1968] = 'd160;
    mem[1969] = 'd160;
    mem[1970] = 'd176;
    mem[1971] = 'd176;
    mem[1972] = 'd220;
    mem[1973] = 'd220;
    mem[1974] = 'd304;
    mem[1975] = 'd308;
    mem[1976] = 'd428;
    mem[1977] = 'd436;
    mem[1978] = 'd628;
    mem[1979] = 'd636;
    mem[1980] = 'd820;
    mem[1981] = 'd840;
    mem[1982] = 'd980;
    mem[1983] = 'd1004;
    mem[1984] = 'd988;
    mem[1985] = 'd1020;
    mem[1986] = 'd984;
    mem[1987] = 'd1020;
    mem[1988] = 'd988;
    mem[1989] = 'd1020;
    mem[1990] = 'd988;
    mem[1991] = 'd1020;
    mem[1992] = 'd944;
    mem[1993] = 'd972;
    mem[1994] = 'd788;
    mem[1995] = 'd804;
    mem[1996] = 'd596;
    mem[1997] = 'd608;
    mem[1998] = 'd408;
    mem[1999] = 'd412;
    mem[2000] = 'd288;
    mem[2001] = 'd296;
    mem[2002] = 'd212;
    mem[2003] = 'd216;
    mem[2004] = 'd172;
    mem[2005] = 'd176;
    mem[2006] = 'd164;
    mem[2007] = 'd160;
    mem[2008] = 'd156;
    mem[2009] = 'd160;
    mem[2010] = 'd168;
    mem[2011] = 'd172;
    mem[2012] = 'd172;
    mem[2013] = 'd176;
    mem[2014] = 'd172;
    mem[2015] = 'd180;
    mem[2016] = 'd168;
    mem[2017] = 'd184;
    mem[2018] = 'd540;
    mem[2019] = 'd860;
    mem[2020] = 'd668;
    mem[2021] = 'd956;
    mem[2022] = 'd1020;
    mem[2023] = 'd1020;
    mem[2024] = 'd1020;
    mem[2025] = 'd1020;
    mem[2026] = 'd1020;
    mem[2027] = 'd1020;
    mem[2028] = 'd1020;
    mem[2029] = 'd1020;
    mem[2030] = 'd936;
    mem[2031] = 'd976;
    mem[2032] = 'd76;
    mem[2033] = 'd564;
    mem[2034] = 'd56;
    mem[2035] = 'd488;
    mem[2036] = 'd88;
    mem[2037] = 'd84;
    mem[2038] = 'd88;
    mem[2039] = 'd88;
    mem[2040] = 'd160;
    mem[2041] = 'd164;
    mem[2042] = 'd432;
    mem[2043] = 'd440;
    mem[2044] = 'd532;
    mem[2045] = 'd544;
    mem[2046] = 'd580;
    mem[2047] = 'd596;
    mem[2048] = 'd596;
    mem[2049] = 'd608;
    mem[2050] = 'd576;
    mem[2051] = 'd588;
    mem[2052] = 'd512;
    mem[2053] = 'd524;
    mem[2054] = 'd412;
    mem[2055] = 'd424;
    mem[2056] = 'd264;
    mem[2057] = 'd268;
    mem[2058] = 'd152;
    mem[2059] = 'd152;
    mem[2060] = 'd192;
    mem[2061] = 'd268;
    mem[2062] = 'd268;
    mem[2063] = 'd508;
    mem[2064] = 'd296;
    mem[2065] = 'd612;
    mem[2066] = 'd284;
    mem[2067] = 'd596;
    mem[2068] = 'd248;
    mem[2069] = 'd472;
    mem[2070] = 'd176;
    mem[2071] = 'd248;
    mem[2072] = 'd180;
    mem[2073] = 'd184;
    mem[2074] = 'd288;
    mem[2075] = 'd292;
    mem[2076] = 'd412;
    mem[2077] = 'd420;
    mem[2078] = 'd488;
    mem[2079] = 'd500;
    mem[2080] = 'd540;
    mem[2081] = 'd548;
    mem[2082] = 'd548;
    mem[2083] = 'd560;
    mem[2084] = 'd528;
    mem[2085] = 'd536;
    mem[2086] = 'd468;
    mem[2087] = 'd480;
    mem[2088] = 'd340;
    mem[2089] = 'd348;
    mem[2090] = 'd116;
    mem[2091] = 'd116;
    mem[2092] = 'd88;
    mem[2093] = 'd88;
    mem[2094] = 'd92;
    mem[2095] = 'd100;
    mem[2096] = 'd44;
    mem[2097] = 'd524;
    mem[2098] = 'd28;
    mem[2099] = 'd536;
    mem[2100] = 'd952;
    mem[2101] = 'd984;
    mem[2102] = 'd1020;
    mem[2103] = 'd1020;
    mem[2104] = 'd1020;
    mem[2105] = 'd1020;
    mem[2106] = 'd1020;
    mem[2107] = 'd1020;
    mem[2108] = 'd976;
    mem[2109] = 'd1000;
    mem[2110] = 'd564;
    mem[2111] = 'd940;
    mem[2112] = 'd488;
    mem[2113] = 'd744;
    mem[2114] = 'd84;
    mem[2115] = 'd84;
    mem[2116] = 'd88;
    mem[2117] = 'd88;
    mem[2118] = 'd164;
    mem[2119] = 'd164;
    mem[2120] = 'd440;
    mem[2121] = 'd432;
    mem[2122] = 'd544;
    mem[2123] = 'd536;
    mem[2124] = 'd596;
    mem[2125] = 'd584;
    mem[2126] = 'd608;
    mem[2127] = 'd600;
    mem[2128] = 'd588;
    mem[2129] = 'd576;
    mem[2130] = 'd524;
    mem[2131] = 'd516;
    mem[2132] = 'd424;
    mem[2133] = 'd416;
    mem[2134] = 'd268;
    mem[2135] = 'd264;
    mem[2136] = 'd152;
    mem[2137] = 'd152;
    mem[2138] = 'd268;
    mem[2139] = 'd272;
    mem[2140] = 'd508;
    mem[2141] = 'd516;
    mem[2142] = 'd612;
    mem[2143] = 'd620;
    mem[2144] = 'd596;
    mem[2145] = 'd604;
    mem[2146] = 'd472;
    mem[2147] = 'd480;
    mem[2148] = 'd248;
    mem[2149] = 'd252;
    mem[2150] = 'd184;
    mem[2151] = 'd184;
    mem[2152] = 'd292;
    mem[2153] = 'd288;
    mem[2154] = 'd420;
    mem[2155] = 'd416;
    mem[2156] = 'd500;
    mem[2157] = 'd492;
    mem[2158] = 'd548;
    mem[2159] = 'd540;
    mem[2160] = 'd560;
    mem[2161] = 'd548;
    mem[2162] = 'd536;
    mem[2163] = 'd528;
    mem[2164] = 'd480;
    mem[2165] = 'd468;
    mem[2166] = 'd348;
    mem[2167] = 'd340;
    mem[2168] = 'd116;
    mem[2169] = 'd116;
    mem[2170] = 'd88;
    mem[2171] = 'd88;
    mem[2172] = 'd100;
    mem[2173] = 'd100;
    mem[2174] = 'd524;
    mem[2175] = 'd796;
    mem[2176] = 'd536;
    mem[2177] = 'd932;
    mem[2178] = 'd984;
    mem[2179] = 'd1004;
    mem[2180] = 'd1020;
    mem[2181] = 'd1020;
    mem[2182] = 'd1020;
    mem[2183] = 'd1020;
    mem[2184] = 'd1020;
    mem[2185] = 'd1020;
    mem[2186] = 'd720;
    mem[2187] = 'd852;
    mem[2188] = 'd16;
    mem[2189] = 'd552;
    mem[2190] = 'd52;
    mem[2191] = 'd632;
    mem[2192] = 'd92;
    mem[2193] = 'd152;
    mem[2194] = 'd84;
    mem[2195] = 'd84;
    mem[2196] = 'd328;
    mem[2197] = 'd332;
    mem[2198] = 'd452;
    mem[2199] = 'd464;
    mem[2200] = 'd508;
    mem[2201] = 'd520;
    mem[2202] = 'd532;
    mem[2203] = 'd544;
    mem[2204] = 'd536;
    mem[2205] = 'd552;
    mem[2206] = 'd540;
    mem[2207] = 'd552;
    mem[2208] = 'd536;
    mem[2209] = 'd548;
    mem[2210] = 'd540;
    mem[2211] = 'd556;
    mem[2212] = 'd564;
    mem[2213] = 'd576;
    mem[2214] = 'd520;
    mem[2215] = 'd532;
    mem[2216] = 'd196;
    mem[2217] = 'd200;
    mem[2218] = 'd100;
    mem[2219] = 'd104;
    mem[2220] = 'd144;
    mem[2221] = 'd144;
    mem[2222] = 'd128;
    mem[2223] = 'd128;
    mem[2224] = 'd100;
    mem[2225] = 'd100;
    mem[2226] = 'd248;
    mem[2227] = 'd252;
    mem[2228] = 'd464;
    mem[2229] = 'd476;
    mem[2230] = 'd480;
    mem[2231] = 'd492;
    mem[2232] = 'd460;
    mem[2233] = 'd472;
    mem[2234] = 'd456;
    mem[2235] = 'd464;
    mem[2236] = 'd452;
    mem[2237] = 'd460;
    mem[2238] = 'd440;
    mem[2239] = 'd452;
    mem[2240] = 'd420;
    mem[2241] = 'd432;
    mem[2242] = 'd388;
    mem[2243] = 'd396;
    mem[2244] = 'd328;
    mem[2245] = 'd336;
    mem[2246] = 'd208;
    mem[2247] = 'd212;
    mem[2248] = 'd84;
    mem[2249] = 'd84;
    mem[2250] = 'd84;
    mem[2251] = 'd212;
    mem[2252] = 'd40;
    mem[2253] = 'd596;
    mem[2254] = 'd12;
    mem[2255] = 'd556;
    mem[2256] = 'd652;
    mem[2257] = 'd816;
    mem[2258] = 'd1020;
    mem[2259] = 'd1020;
    mem[2260] = 'd1020;
    mem[2261] = 'd1020;
    mem[2262] = 'd1020;
    mem[2263] = 'd1020;
    mem[2264] = 'd852;
    mem[2265] = 'd972;
    mem[2266] = 'd552;
    mem[2267] = 'd948;
    mem[2268] = 'd632;
    mem[2269] = 'd952;
    mem[2270] = 'd152;
    mem[2271] = 'd184;
    mem[2272] = 'd84;
    mem[2273] = 'd84;
    mem[2274] = 'd332;
    mem[2275] = 'd328;
    mem[2276] = 'd464;
    mem[2277] = 'd452;
    mem[2278] = 'd520;
    mem[2279] = 'd512;
    mem[2280] = 'd544;
    mem[2281] = 'd536;
    mem[2282] = 'd552;
    mem[2283] = 'd540;
    mem[2284] = 'd552;
    mem[2285] = 'd540;
    mem[2286] = 'd548;
    mem[2287] = 'd540;
    mem[2288] = 'd556;
    mem[2289] = 'd544;
    mem[2290] = 'd576;
    mem[2291] = 'd564;
    mem[2292] = 'd532;
    mem[2293] = 'd520;
    mem[2294] = 'd200;
    mem[2295] = 'd196;
    mem[2296] = 'd104;
    mem[2297] = 'd100;
    mem[2298] = 'd144;
    mem[2299] = 'd144;
    mem[2300] = 'd128;
    mem[2301] = 'd128;
    mem[2302] = 'd100;
    mem[2303] = 'd100;
    mem[2304] = 'd252;
    mem[2305] = 'd248;
    mem[2306] = 'd476;
    mem[2307] = 'd464;
    mem[2308] = 'd492;
    mem[2309] = 'd484;
    mem[2310] = 'd472;
    mem[2311] = 'd460;
    mem[2312] = 'd464;
    mem[2313] = 'd456;
    mem[2314] = 'd460;
    mem[2315] = 'd452;
    mem[2316] = 'd452;
    mem[2317] = 'd444;
    mem[2318] = 'd432;
    mem[2319] = 'd424;
    mem[2320] = 'd396;
    mem[2321] = 'd388;
    mem[2322] = 'd336;
    mem[2323] = 'd332;
    mem[2324] = 'd212;
    mem[2325] = 'd208;
    mem[2326] = 'd84;
    mem[2327] = 'd84;
    mem[2328] = 'd212;
    mem[2329] = 'd280;
    mem[2330] = 'd596;
    mem[2331] = 'd896;
    mem[2332] = 'd556;
    mem[2333] = 'd932;
    mem[2334] = 'd816;
    mem[2335] = 'd960;
    mem[2336] = 'd1020;
    mem[2337] = 'd1020;
    mem[2338] = 'd1020;
    mem[2339] = 'd1020;
    mem[2340] = 'd1020;
    mem[2341] = 'd1020;
    mem[2342] = 'd464;
    mem[2343] = 'd716;
    mem[2344] = 'd20;
    mem[2345] = 'd572;
    mem[2346] = 'd72;
    mem[2347] = 'd640;
    mem[2348] = 'd96;
    mem[2349] = 'd384;
    mem[2350] = 'd92;
    mem[2351] = 'd88;
    mem[2352] = 'd212;
    mem[2353] = 'd216;
    mem[2354] = 'd252;
    mem[2355] = 'd256;
    mem[2356] = 'd260;
    mem[2357] = 'd268;
    mem[2358] = 'd272;
    mem[2359] = 'd280;
    mem[2360] = 'd280;
    mem[2361] = 'd292;
    mem[2362] = 'd280;
    mem[2363] = 'd288;
    mem[2364] = 'd264;
    mem[2365] = 'd268;
    mem[2366] = 'd244;
    mem[2367] = 'd252;
    mem[2368] = 'd232;
    mem[2369] = 'd236;
    mem[2370] = 'd216;
    mem[2371] = 'd224;
    mem[2372] = 'd144;
    mem[2373] = 'd148;
    mem[2374] = 'd84;
    mem[2375] = 'd84;
    mem[2376] = 'd76;
    mem[2377] = 'd264;
    mem[2378] = 'd76;
    mem[2379] = 'd188;
    mem[2380] = 'd84;
    mem[2381] = 'd84;
    mem[2382] = 'd148;
    mem[2383] = 'd152;
    mem[2384] = 'd180;
    mem[2385] = 'd184;
    mem[2386] = 'd180;
    mem[2387] = 'd188;
    mem[2388] = 'd184;
    mem[2389] = 'd188;
    mem[2390] = 'd192;
    mem[2391] = 'd196;
    mem[2392] = 'd196;
    mem[2393] = 'd200;
    mem[2394] = 'd184;
    mem[2395] = 'd188;
    mem[2396] = 'd168;
    mem[2397] = 'd172;
    mem[2398] = 'd148;
    mem[2399] = 'd156;
    mem[2400] = 'd136;
    mem[2401] = 'd140;
    mem[2402] = 'd104;
    mem[2403] = 'd104;
    mem[2404] = 'd92;
    mem[2405] = 'd88;
    mem[2406] = 'd68;
    mem[2407] = 'd420;
    mem[2408] = 'd56;
    mem[2409] = 'd612;
    mem[2410] = 'd20;
    mem[2411] = 'd572;
    mem[2412] = 'd420;
    mem[2413] = 'd692;
    mem[2414] = 'd1020;
    mem[2415] = 'd1020;
    mem[2416] = 'd1020;
    mem[2417] = 'd1020;
    mem[2418] = 'd1020;
    mem[2419] = 'd1020;
    mem[2420] = 'd716;
    mem[2421] = 'd940;
    mem[2422] = 'd572;
    mem[2423] = 'd956;
    mem[2424] = 'd640;
    mem[2425] = 'd948;
    mem[2426] = 'd384;
    mem[2427] = 'd524;
    mem[2428] = 'd88;
    mem[2429] = 'd88;
    mem[2430] = 'd216;
    mem[2431] = 'd212;
    mem[2432] = 'd256;
    mem[2433] = 'd252;
    mem[2434] = 'd268;
    mem[2435] = 'd264;
    mem[2436] = 'd280;
    mem[2437] = 'd276;
    mem[2438] = 'd292;
    mem[2439] = 'd284;
    mem[2440] = 'd288;
    mem[2441] = 'd280;
    mem[2442] = 'd268;
    mem[2443] = 'd264;
    mem[2444] = 'd252;
    mem[2445] = 'd244;
    mem[2446] = 'd236;
    mem[2447] = 'd232;
    mem[2448] = 'd224;
    mem[2449] = 'd220;
    mem[2450] = 'd148;
    mem[2451] = 'd144;
    mem[2452] = 'd84;
    mem[2453] = 'd84;
    mem[2454] = 'd264;
    mem[2455] = 'd320;
    mem[2456] = 'd188;
    mem[2457] = 'd220;
    mem[2458] = 'd84;
    mem[2459] = 'd84;
    mem[2460] = 'd152;
    mem[2461] = 'd148;
    mem[2462] = 'd184;
    mem[2463] = 'd180;
    mem[2464] = 'd188;
    mem[2465] = 'd180;
    mem[2466] = 'd188;
    mem[2467] = 'd188;
    mem[2468] = 'd196;
    mem[2469] = 'd192;
    mem[2470] = 'd200;
    mem[2471] = 'd196;
    mem[2472] = 'd188;
    mem[2473] = 'd184;
    mem[2474] = 'd172;
    mem[2475] = 'd168;
    mem[2476] = 'd156;
    mem[2477] = 'd148;
    mem[2478] = 'd140;
    mem[2479] = 'd140;
    mem[2480] = 'd104;
    mem[2481] = 'd104;
    mem[2482] = 'd88;
    mem[2483] = 'd88;
    mem[2484] = 'd420;
    mem[2485] = 'd600;
    mem[2486] = 'd612;
    mem[2487] = 'd908;
    mem[2488] = 'd572;
    mem[2489] = 'd948;
    mem[2490] = 'd692;
    mem[2491] = 'd940;
    mem[2492] = 'd1020;
    mem[2493] = 'd1020;
    mem[2494] = 'd1020;
    mem[2495] = 'd1020;
    mem[2496] = 'd1020;
    mem[2497] = 'd1020;
    mem[2498] = 'd288;
    mem[2499] = 'd616;
    mem[2500] = 'd24;
    mem[2501] = 'd588;
    mem[2502] = 'd76;
    mem[2503] = 'd652;
    mem[2504] = 'd84;
    mem[2505] = 'd540;
    mem[2506] = 'd92;
    mem[2507] = 'd96;
    mem[2508] = 'd88;
    mem[2509] = 'd88;
    mem[2510] = 'd104;
    mem[2511] = 'd104;
    mem[2512] = 'd112;
    mem[2513] = 'd116;
    mem[2514] = 'd124;
    mem[2515] = 'd128;
    mem[2516] = 'd136;
    mem[2517] = 'd144;
    mem[2518] = 'd148;
    mem[2519] = 'd156;
    mem[2520] = 'd148;
    mem[2521] = 'd152;
    mem[2522] = 'd144;
    mem[2523] = 'd148;
    mem[2524] = 'd148;
    mem[2525] = 'd152;
    mem[2526] = 'd128;
    mem[2527] = 'd132;
    mem[2528] = 'd108;
    mem[2529] = 'd108;
    mem[2530] = 'd80;
    mem[2531] = 'd80;
    mem[2532] = 'd136;
    mem[2533] = 'd704;
    mem[2534] = 'd124;
    mem[2535] = 'd568;
    mem[2536] = 'd84;
    mem[2537] = 'd84;
    mem[2538] = 'd116;
    mem[2539] = 'd120;
    mem[2540] = 'd160;
    mem[2541] = 'd168;
    mem[2542] = 'd176;
    mem[2543] = 'd180;
    mem[2544] = 'd180;
    mem[2545] = 'd184;
    mem[2546] = 'd192;
    mem[2547] = 'd196;
    mem[2548] = 'd196;
    mem[2549] = 'd204;
    mem[2550] = 'd188;
    mem[2551] = 'd196;
    mem[2552] = 'd180;
    mem[2553] = 'd184;
    mem[2554] = 'd172;
    mem[2555] = 'd176;
    mem[2556] = 'd160;
    mem[2557] = 'd160;
    mem[2558] = 'd124;
    mem[2559] = 'd128;
    mem[2560] = 'd96;
    mem[2561] = 'd108;
    mem[2562] = 'd44;
    mem[2563] = 'd552;
    mem[2564] = 'd68;
    mem[2565] = 'd636;
    mem[2566] = 'd28;
    mem[2567] = 'd588;
    mem[2568] = 'd240;
    mem[2569] = 'd600;
    mem[2570] = 'd1020;
    mem[2571] = 'd1020;
    mem[2572] = 'd1020;
    mem[2573] = 'd1020;
    mem[2574] = 'd1020;
    mem[2575] = 'd1020;
    mem[2576] = 'd616;
    mem[2577] = 'd920;
    mem[2578] = 'd588;
    mem[2579] = 'd956;
    mem[2580] = 'd652;
    mem[2581] = 'd960;
    mem[2582] = 'd540;
    mem[2583] = 'd768;
    mem[2584] = 'd96;
    mem[2585] = 'd96;
    mem[2586] = 'd88;
    mem[2587] = 'd88;
    mem[2588] = 'd104;
    mem[2589] = 'd104;
    mem[2590] = 'd116;
    mem[2591] = 'd112;
    mem[2592] = 'd128;
    mem[2593] = 'd124;
    mem[2594] = 'd144;
    mem[2595] = 'd140;
    mem[2596] = 'd156;
    mem[2597] = 'd148;
    mem[2598] = 'd152;
    mem[2599] = 'd148;
    mem[2600] = 'd148;
    mem[2601] = 'd144;
    mem[2602] = 'd152;
    mem[2603] = 'd148;
    mem[2604] = 'd132;
    mem[2605] = 'd128;
    mem[2606] = 'd108;
    mem[2607] = 'd108;
    mem[2608] = 'd80;
    mem[2609] = 'd76;
    mem[2610] = 'd704;
    mem[2611] = 'd844;
    mem[2612] = 'd568;
    mem[2613] = 'd672;
    mem[2614] = 'd84;
    mem[2615] = 'd80;
    mem[2616] = 'd120;
    mem[2617] = 'd120;
    mem[2618] = 'd168;
    mem[2619] = 'd164;
    mem[2620] = 'd180;
    mem[2621] = 'd172;
    mem[2622] = 'd184;
    mem[2623] = 'd180;
    mem[2624] = 'd196;
    mem[2625] = 'd192;
    mem[2626] = 'd204;
    mem[2627] = 'd200;
    mem[2628] = 'd196;
    mem[2629] = 'd192;
    mem[2630] = 'd184;
    mem[2631] = 'd180;
    mem[2632] = 'd176;
    mem[2633] = 'd172;
    mem[2634] = 'd160;
    mem[2635] = 'd160;
    mem[2636] = 'd128;
    mem[2637] = 'd124;
    mem[2638] = 'd108;
    mem[2639] = 'd112;
    mem[2640] = 'd552;
    mem[2641] = 'd812;
    mem[2642] = 'd636;
    mem[2643] = 'd936;
    mem[2644] = 'd588;
    mem[2645] = 'd960;
    mem[2646] = 'd600;
    mem[2647] = 'd912;
    mem[2648] = 'd1020;
    mem[2649] = 'd1020;
    mem[2650] = 'd1020;
    mem[2651] = 'd1020;
    mem[2652] = 'd1020;
    mem[2653] = 'd1020;
    mem[2654] = 'd168;
    mem[2655] = 'd556;
    mem[2656] = 'd28;
    mem[2657] = 'd588;
    mem[2658] = 'd68;
    mem[2659] = 'd660;
    mem[2660] = 'd68;
    mem[2661] = 'd624;
    mem[2662] = 'd88;
    mem[2663] = 'd192;
    mem[2664] = 'd108;
    mem[2665] = 'd108;
    mem[2666] = 'd132;
    mem[2667] = 'd136;
    mem[2668] = 'd164;
    mem[2669] = 'd168;
    mem[2670] = 'd176;
    mem[2671] = 'd180;
    mem[2672] = 'd180;
    mem[2673] = 'd184;
    mem[2674] = 'd180;
    mem[2675] = 'd184;
    mem[2676] = 'd184;
    mem[2677] = 'd192;
    mem[2678] = 'd188;
    mem[2679] = 'd196;
    mem[2680] = 'd180;
    mem[2681] = 'd184;
    mem[2682] = 'd128;
    mem[2683] = 'd132;
    mem[2684] = 'd116;
    mem[2685] = 'd120;
    mem[2686] = 'd88;
    mem[2687] = 'd260;
    mem[2688] = 'd180;
    mem[2689] = 'd876;
    mem[2690] = 'd168;
    mem[2691] = 'd848;
    mem[2692] = 'd80;
    mem[2693] = 'd156;
    mem[2694] = 'd120;
    mem[2695] = 'd120;
    mem[2696] = 'd172;
    mem[2697] = 'd176;
    mem[2698] = 'd208;
    mem[2699] = 'd212;
    mem[2700] = 'd212;
    mem[2701] = 'd216;
    mem[2702] = 'd208;
    mem[2703] = 'd212;
    mem[2704] = 'd204;
    mem[2705] = 'd212;
    mem[2706] = 'd212;
    mem[2707] = 'd216;
    mem[2708] = 'd212;
    mem[2709] = 'd216;
    mem[2710] = 'd200;
    mem[2711] = 'd204;
    mem[2712] = 'd160;
    mem[2713] = 'd164;
    mem[2714] = 'd136;
    mem[2715] = 'd136;
    mem[2716] = 'd76;
    mem[2717] = 'd224;
    mem[2718] = 'd40;
    mem[2719] = 'd596;
    mem[2720] = 'd68;
    mem[2721] = 'd652;
    mem[2722] = 'd32;
    mem[2723] = 'd592;
    mem[2724] = 'd136;
    mem[2725] = 'd540;
    mem[2726] = 'd1020;
    mem[2727] = 'd1020;
    mem[2728] = 'd1020;
    mem[2729] = 'd1020;
    mem[2730] = 'd1020;
    mem[2731] = 'd1020;
    mem[2732] = 'd556;
    mem[2733] = 'd896;
    mem[2734] = 'd588;
    mem[2735] = 'd956;
    mem[2736] = 'd660;
    mem[2737] = 'd972;
    mem[2738] = 'd624;
    mem[2739] = 'd904;
    mem[2740] = 'd192;
    mem[2741] = 'd240;
    mem[2742] = 'd108;
    mem[2743] = 'd108;
    mem[2744] = 'd136;
    mem[2745] = 'd132;
    mem[2746] = 'd168;
    mem[2747] = 'd164;
    mem[2748] = 'd180;
    mem[2749] = 'd176;
    mem[2750] = 'd184;
    mem[2751] = 'd180;
    mem[2752] = 'd184;
    mem[2753] = 'd180;
    mem[2754] = 'd192;
    mem[2755] = 'd188;
    mem[2756] = 'd196;
    mem[2757] = 'd192;
    mem[2758] = 'd184;
    mem[2759] = 'd180;
    mem[2760] = 'd132;
    mem[2761] = 'd128;
    mem[2762] = 'd120;
    mem[2763] = 'd116;
    mem[2764] = 'd260;
    mem[2765] = 'd296;
    mem[2766] = 'd876;
    mem[2767] = 'd1004;
    mem[2768] = 'd848;
    mem[2769] = 'd980;
    mem[2770] = 'd156;
    mem[2771] = 'd176;
    mem[2772] = 'd120;
    mem[2773] = 'd120;
    mem[2774] = 'd176;
    mem[2775] = 'd172;
    mem[2776] = 'd212;
    mem[2777] = 'd208;
    mem[2778] = 'd216;
    mem[2779] = 'd212;
    mem[2780] = 'd212;
    mem[2781] = 'd208;
    mem[2782] = 'd212;
    mem[2783] = 'd204;
    mem[2784] = 'd216;
    mem[2785] = 'd212;
    mem[2786] = 'd216;
    mem[2787] = 'd216;
    mem[2788] = 'd204;
    mem[2789] = 'd200;
    mem[2790] = 'd164;
    mem[2791] = 'd160;
    mem[2792] = 'd136;
    mem[2793] = 'd136;
    mem[2794] = 'd224;
    mem[2795] = 'd304;
    mem[2796] = 'd596;
    mem[2797] = 'd880;
    mem[2798] = 'd652;
    mem[2799] = 'd960;
    mem[2800] = 'd592;
    mem[2801] = 'd956;
    mem[2802] = 'd540;
    mem[2803] = 'd892;
    mem[2804] = 'd1020;
    mem[2805] = 'd1020;
    mem[2806] = 'd1020;
    mem[2807] = 'd1020;
    mem[2808] = 'd1020;
    mem[2809] = 'd1020;
    mem[2810] = 'd124;
    mem[2811] = 'd528;
    mem[2812] = 'd28;
    mem[2813] = 'd584;
    mem[2814] = 'd60;
    mem[2815] = 'd664;
    mem[2816] = 'd72;
    mem[2817] = 'd648;
    mem[2818] = 'd76;
    mem[2819] = 'd408;
    mem[2820] = 'd120;
    mem[2821] = 'd120;
    mem[2822] = 'd120;
    mem[2823] = 'd124;
    mem[2824] = 'd168;
    mem[2825] = 'd168;
    mem[2826] = 'd188;
    mem[2827] = 'd188;
    mem[2828] = 'd192;
    mem[2829] = 'd192;
    mem[2830] = 'd192;
    mem[2831] = 'd196;
    mem[2832] = 'd192;
    mem[2833] = 'd200;
    mem[2834] = 'd188;
    mem[2835] = 'd188;
    mem[2836] = 'd140;
    mem[2837] = 'd144;
    mem[2838] = 'd124;
    mem[2839] = 'd124;
    mem[2840] = 'd88;
    mem[2841] = 'd84;
    mem[2842] = 'd136;
    mem[2843] = 'd644;
    mem[2844] = 'd192;
    mem[2845] = 'd888;
    mem[2846] = 'd188;
    mem[2847] = 'd880;
    mem[2848] = 'd120;
    mem[2849] = 'd540;
    mem[2850] = 'd100;
    mem[2851] = 'd96;
    mem[2852] = 'd128;
    mem[2853] = 'd132;
    mem[2854] = 'd176;
    mem[2855] = 'd180;
    mem[2856] = 'd204;
    mem[2857] = 'd208;
    mem[2858] = 'd204;
    mem[2859] = 'd208;
    mem[2860] = 'd200;
    mem[2861] = 'd208;
    mem[2862] = 'd204;
    mem[2863] = 'd208;
    mem[2864] = 'd204;
    mem[2865] = 'd208;
    mem[2866] = 'd176;
    mem[2867] = 'd180;
    mem[2868] = 'd116;
    mem[2869] = 'd120;
    mem[2870] = 'd120;
    mem[2871] = 'd116;
    mem[2872] = 'd48;
    mem[2873] = 'd444;
    mem[2874] = 'd56;
    mem[2875] = 'd620;
    mem[2876] = 'd64;
    mem[2877] = 'd664;
    mem[2878] = 'd28;
    mem[2879] = 'd588;
    mem[2880] = 'd88;
    mem[2881] = 'd512;
    mem[2882] = 'd1012;
    mem[2883] = 'd1012;
    mem[2884] = 'd1020;
    mem[2885] = 'd1020;
    mem[2886] = 'd1020;
    mem[2887] = 'd1020;
    mem[2888] = 'd528;
    mem[2889] = 'd880;
    mem[2890] = 'd584;
    mem[2891] = 'd948;
    mem[2892] = 'd664;
    mem[2893] = 'd980;
    mem[2894] = 'd648;
    mem[2895] = 'd940;
    mem[2896] = 'd408;
    mem[2897] = 'd572;
    mem[2898] = 'd120;
    mem[2899] = 'd120;
    mem[2900] = 'd124;
    mem[2901] = 'd120;
    mem[2902] = 'd168;
    mem[2903] = 'd168;
    mem[2904] = 'd188;
    mem[2905] = 'd188;
    mem[2906] = 'd192;
    mem[2907] = 'd192;
    mem[2908] = 'd196;
    mem[2909] = 'd192;
    mem[2910] = 'd200;
    mem[2911] = 'd196;
    mem[2912] = 'd188;
    mem[2913] = 'd188;
    mem[2914] = 'd144;
    mem[2915] = 'd140;
    mem[2916] = 'd124;
    mem[2917] = 'd124;
    mem[2918] = 'd84;
    mem[2919] = 'd84;
    mem[2920] = 'd644;
    mem[2921] = 'd752;
    mem[2922] = 'd888;
    mem[2923] = 'd1016;
    mem[2924] = 'd880;
    mem[2925] = 'd1012;
    mem[2926] = 'd540;
    mem[2927] = 'd636;
    mem[2928] = 'd96;
    mem[2929] = 'd96;
    mem[2930] = 'd132;
    mem[2931] = 'd128;
    mem[2932] = 'd180;
    mem[2933] = 'd176;
    mem[2934] = 'd208;
    mem[2935] = 'd204;
    mem[2936] = 'd208;
    mem[2937] = 'd208;
    mem[2938] = 'd208;
    mem[2939] = 'd204;
    mem[2940] = 'd208;
    mem[2941] = 'd208;
    mem[2942] = 'd208;
    mem[2943] = 'd204;
    mem[2944] = 'd180;
    mem[2945] = 'd176;
    mem[2946] = 'd120;
    mem[2947] = 'd116;
    mem[2948] = 'd116;
    mem[2949] = 'd112;
    mem[2950] = 'd444;
    mem[2951] = 'd648;
    mem[2952] = 'd620;
    mem[2953] = 'd904;
    mem[2954] = 'd664;
    mem[2955] = 'd980;
    mem[2956] = 'd588;
    mem[2957] = 'd948;
    mem[2958] = 'd512;
    mem[2959] = 'd876;
    mem[2960] = 'd1012;
    mem[2961] = 'd1016;
    mem[2962] = 'd1020;
    mem[2963] = 'd1020;
    mem[2964] = 'd1020;
    mem[2965] = 'd1020;
    mem[2966] = 'd120;
    mem[2967] = 'd520;
    mem[2968] = 'd28;
    mem[2969] = 'd576;
    mem[2970] = 'd56;
    mem[2971] = 'd660;
    mem[2972] = 'd92;
    mem[2973] = 'd684;
    mem[2974] = 'd72;
    mem[2975] = 'd608;
    mem[2976] = 'd92;
    mem[2977] = 'd200;
    mem[2978] = 'd128;
    mem[2979] = 'd132;
    mem[2980] = 'd108;
    mem[2981] = 'd112;
    mem[2982] = 'd120;
    mem[2983] = 'd124;
    mem[2984] = 'd136;
    mem[2985] = 'd140;
    mem[2986] = 'd144;
    mem[2987] = 'd148;
    mem[2988] = 'd140;
    mem[2989] = 'd140;
    mem[2990] = 'd112;
    mem[2991] = 'd116;
    mem[2992] = 'd112;
    mem[2993] = 'd116;
    mem[2994] = 'd104;
    mem[2995] = 'd104;
    mem[2996] = 'd92;
    mem[2997] = 'd356;
    mem[2998] = 'd176;
    mem[2999] = 'd856;
    mem[3000] = 'd196;
    mem[3001] = 'd884;
    mem[3002] = 'd192;
    mem[3003] = 'd884;
    mem[3004] = 'd172;
    mem[3005] = 'd840;
    mem[3006] = 'd80;
    mem[3007] = 'd268;
    mem[3008] = 'd120;
    mem[3009] = 'd120;
    mem[3010] = 'd120;
    mem[3011] = 'd120;
    mem[3012] = 'd120;
    mem[3013] = 'd124;
    mem[3014] = 'd128;
    mem[3015] = 'd132;
    mem[3016] = 'd132;
    mem[3017] = 'd136;
    mem[3018] = 'd136;
    mem[3019] = 'd136;
    mem[3020] = 'd124;
    mem[3021] = 'd128;
    mem[3022] = 'd100;
    mem[3023] = 'd100;
    mem[3024] = 'd124;
    mem[3025] = 'd128;
    mem[3026] = 'd68;
    mem[3027] = 'd220;
    mem[3028] = 'd40;
    mem[3029] = 'd588;
    mem[3030] = 'd84;
    mem[3031] = 'd668;
    mem[3032] = 'd60;
    mem[3033] = 'd668;
    mem[3034] = 'd28;
    mem[3035] = 'd580;
    mem[3036] = 'd88;
    mem[3037] = 'd504;
    mem[3038] = 'd1012;
    mem[3039] = 'd1012;
    mem[3040] = 'd1020;
    mem[3041] = 'd1020;
    mem[3042] = 'd1020;
    mem[3043] = 'd1020;
    mem[3044] = 'd520;
    mem[3045] = 'd872;
    mem[3046] = 'd576;
    mem[3047] = 'd932;
    mem[3048] = 'd660;
    mem[3049] = 'd984;
    mem[3050] = 'd684;
    mem[3051] = 'd968;
    mem[3052] = 'd608;
    mem[3053] = 'd876;
    mem[3054] = 'd200;
    mem[3055] = 'd256;
    mem[3056] = 'd132;
    mem[3057] = 'd128;
    mem[3058] = 'd112;
    mem[3059] = 'd112;
    mem[3060] = 'd124;
    mem[3061] = 'd120;
    mem[3062] = 'd140;
    mem[3063] = 'd140;
    mem[3064] = 'd148;
    mem[3065] = 'd144;
    mem[3066] = 'd140;
    mem[3067] = 'd140;
    mem[3068] = 'd116;
    mem[3069] = 'd112;
    mem[3070] = 'd116;
    mem[3071] = 'd112;
    mem[3072] = 'd104;
    mem[3073] = 'd100;
    mem[3074] = 'd356;
    mem[3075] = 'd432;
    mem[3076] = 'd856;
    mem[3077] = 'd1008;
    mem[3078] = 'd884;
    mem[3079] = 'd1020;
    mem[3080] = 'd884;
    mem[3081] = 'd1020;
    mem[3082] = 'd840;
    mem[3083] = 'd992;
    mem[3084] = 'd268;
    mem[3085] = 'd324;
    mem[3086] = 'd120;
    mem[3087] = 'd120;
    mem[3088] = 'd120;
    mem[3089] = 'd120;
    mem[3090] = 'd124;
    mem[3091] = 'd120;
    mem[3092] = 'd132;
    mem[3093] = 'd132;
    mem[3094] = 'd136;
    mem[3095] = 'd136;
    mem[3096] = 'd136;
    mem[3097] = 'd132;
    mem[3098] = 'd128;
    mem[3099] = 'd124;
    mem[3100] = 'd100;
    mem[3101] = 'd100;
    mem[3102] = 'd128;
    mem[3103] = 'd128;
    mem[3104] = 'd220;
    mem[3105] = 'd300;
    mem[3106] = 'd588;
    mem[3107] = 'd872;
    mem[3108] = 'd668;
    mem[3109] = 'd956;
    mem[3110] = 'd668;
    mem[3111] = 'd984;
    mem[3112] = 'd580;
    mem[3113] = 'd940;
    mem[3114] = 'd504;
    mem[3115] = 'd872;
    mem[3116] = 'd1012;
    mem[3117] = 'd1016;
    mem[3118] = 'd1020;
    mem[3119] = 'd1020;
    mem[3120] = 'd1020;
    mem[3121] = 'd1020;
    mem[3122] = 'd168;
    mem[3123] = 'd536;
    mem[3124] = 'd24;
    mem[3125] = 'd560;
    mem[3126] = 'd48;
    mem[3127] = 'd648;
    mem[3128] = 'd104;
    mem[3129] = 'd700;
    mem[3130] = 'd112;
    mem[3131] = 'd680;
    mem[3132] = 'd76;
    mem[3133] = 'd548;
    mem[3134] = 'd84;
    mem[3135] = 'd168;
    mem[3136] = 'd132;
    mem[3137] = 'd132;
    mem[3138] = 'd152;
    mem[3139] = 'd152;
    mem[3140] = 'd152;
    mem[3141] = 'd152;
    mem[3142] = 'd152;
    mem[3143] = 'd156;
    mem[3144] = 'd144;
    mem[3145] = 'd144;
    mem[3146] = 'd136;
    mem[3147] = 'd136;
    mem[3148] = 'd88;
    mem[3149] = 'd88;
    mem[3150] = 'd84;
    mem[3151] = 'd360;
    mem[3152] = 'd164;
    mem[3153] = 'd816;
    mem[3154] = 'd196;
    mem[3155] = 'd868;
    mem[3156] = 'd200;
    mem[3157] = 'd876;
    mem[3158] = 'd196;
    mem[3159] = 'd876;
    mem[3160] = 'd196;
    mem[3161] = 'd868;
    mem[3162] = 'd152;
    mem[3163] = 'd780;
    mem[3164] = 'd76;
    mem[3165] = 'd288;
    mem[3166] = 'd104;
    mem[3167] = 'd100;
    mem[3168] = 'd156;
    mem[3169] = 'd156;
    mem[3170] = 'd152;
    mem[3171] = 'd152;
    mem[3172] = 'd148;
    mem[3173] = 'd152;
    mem[3174] = 'd144;
    mem[3175] = 'd148;
    mem[3176] = 'd140;
    mem[3177] = 'd144;
    mem[3178] = 'd132;
    mem[3179] = 'd128;
    mem[3180] = 'd68;
    mem[3181] = 'd164;
    mem[3182] = 'd44;
    mem[3183] = 'd556;
    mem[3184] = 'd96;
    mem[3185] = 'd660;
    mem[3186] = 'd100;
    mem[3187] = 'd700;
    mem[3188] = 'd52;
    mem[3189] = 'd652;
    mem[3190] = 'd28;
    mem[3191] = 'd568;
    mem[3192] = 'd136;
    mem[3193] = 'd520;
    mem[3194] = 'd1020;
    mem[3195] = 'd1020;
    mem[3196] = 'd1020;
    mem[3197] = 'd1020;
    mem[3198] = 'd1020;
    mem[3199] = 'd1020;
    mem[3200] = 'd536;
    mem[3201] = 'd868;
    mem[3202] = 'd560;
    mem[3203] = 'd924;
    mem[3204] = 'd648;
    mem[3205] = 'd976;
    mem[3206] = 'd700;
    mem[3207] = 'd996;
    mem[3208] = 'd680;
    mem[3209] = 'd956;
    mem[3210] = 'd548;
    mem[3211] = 'd780;
    mem[3212] = 'd168;
    mem[3213] = 'd208;
    mem[3214] = 'd132;
    mem[3215] = 'd128;
    mem[3216] = 'd152;
    mem[3217] = 'd152;
    mem[3218] = 'd152;
    mem[3219] = 'd152;
    mem[3220] = 'd156;
    mem[3221] = 'd152;
    mem[3222] = 'd144;
    mem[3223] = 'd144;
    mem[3224] = 'd136;
    mem[3225] = 'd136;
    mem[3226] = 'd88;
    mem[3227] = 'd88;
    mem[3228] = 'd360;
    mem[3229] = 'd452;
    mem[3230] = 'd816;
    mem[3231] = 'd984;
    mem[3232] = 'd868;
    mem[3233] = 'd1016;
    mem[3234] = 'd876;
    mem[3235] = 'd1020;
    mem[3236] = 'd876;
    mem[3237] = 'd1020;
    mem[3238] = 'd868;
    mem[3239] = 'd1016;
    mem[3240] = 'd780;
    mem[3241] = 'd956;
    mem[3242] = 'd288;
    mem[3243] = 'd356;
    mem[3244] = 'd100;
    mem[3245] = 'd100;
    mem[3246] = 'd156;
    mem[3247] = 'd156;
    mem[3248] = 'd152;
    mem[3249] = 'd152;
    mem[3250] = 'd152;
    mem[3251] = 'd148;
    mem[3252] = 'd148;
    mem[3253] = 'd144;
    mem[3254] = 'd144;
    mem[3255] = 'd140;
    mem[3256] = 'd128;
    mem[3257] = 'd124;
    mem[3258] = 'd164;
    mem[3259] = 'd216;
    mem[3260] = 'd556;
    mem[3261] = 'd816;
    mem[3262] = 'd660;
    mem[3263] = 'd936;
    mem[3264] = 'd700;
    mem[3265] = 'd996;
    mem[3266] = 'd652;
    mem[3267] = 'd980;
    mem[3268] = 'd568;
    mem[3269] = 'd928;
    mem[3270] = 'd520;
    mem[3271] = 'd864;
    mem[3272] = 'd1020;
    mem[3273] = 'd1020;
    mem[3274] = 'd1020;
    mem[3275] = 'd1020;
    mem[3276] = 'd1020;
    mem[3277] = 'd1020;
    mem[3278] = 'd280;
    mem[3279] = 'd592;
    mem[3280] = 'd24;
    mem[3281] = 'd540;
    mem[3282] = 'd44;
    mem[3283] = 'd632;
    mem[3284] = 'd88;
    mem[3285] = 'd700;
    mem[3286] = 'd140;
    mem[3287] = 'd728;
    mem[3288] = 'd144;
    mem[3289] = 'd708;
    mem[3290] = 'd108;
    mem[3291] = 'd640;
    mem[3292] = 'd84;
    mem[3293] = 'd440;
    mem[3294] = 'd76;
    mem[3295] = 'd268;
    mem[3296] = 'd72;
    mem[3297] = 'd184;
    mem[3298] = 'd72;
    mem[3299] = 'd156;
    mem[3300] = 'd72;
    mem[3301] = 'd204;
    mem[3302] = 'd88;
    mem[3303] = 'd336;
    mem[3304] = 'd132;
    mem[3305] = 'd636;
    mem[3306] = 'd184;
    mem[3307] = 'd828;
    mem[3308] = 'd208;
    mem[3309] = 'd856;
    mem[3310] = 'd208;
    mem[3311] = 'd864;
    mem[3312] = 'd204;
    mem[3313] = 'd864;
    mem[3314] = 'd208;
    mem[3315] = 'd864;
    mem[3316] = 'd208;
    mem[3317] = 'd864;
    mem[3318] = 'd204;
    mem[3319] = 'd856;
    mem[3320] = 'd176;
    mem[3321] = 'd812;
    mem[3322] = 'd108;
    mem[3323] = 'd572;
    mem[3324] = 'd72;
    mem[3325] = 'd292;
    mem[3326] = 'd64;
    mem[3327] = 'd188;
    mem[3328] = 'd64;
    mem[3329] = 'd148;
    mem[3330] = 'd64;
    mem[3331] = 'd176;
    mem[3332] = 'd60;
    mem[3333] = 'd276;
    mem[3334] = 'd60;
    mem[3335] = 'd428;
    mem[3336] = 'd76;
    mem[3337] = 'd632;
    mem[3338] = 'd132;
    mem[3339] = 'd692;
    mem[3340] = 'd140;
    mem[3341] = 'd724;
    mem[3342] = 'd84;
    mem[3343] = 'd700;
    mem[3344] = 'd48;
    mem[3345] = 'd636;
    mem[3346] = 'd28;
    mem[3347] = 'd548;
    mem[3348] = 'd236;
    mem[3349] = 'd568;
    mem[3350] = 'd1020;
    mem[3351] = 'd1020;
    mem[3352] = 'd1020;
    mem[3353] = 'd1020;
    mem[3354] = 'd1020;
    mem[3355] = 'd1020;
    mem[3356] = 'd592;
    mem[3357] = 'd876;
    mem[3358] = 'd540;
    mem[3359] = 'd908;
    mem[3360] = 'd632;
    mem[3361] = 'd960;
    mem[3362] = 'd700;
    mem[3363] = 'd1000;
    mem[3364] = 'd728;
    mem[3365] = 'd1004;
    mem[3366] = 'd708;
    mem[3367] = 'd976;
    mem[3368] = 'd640;
    mem[3369] = 'd888;
    mem[3370] = 'd440;
    mem[3371] = 'd604;
    mem[3372] = 'd268;
    mem[3373] = 'd360;
    mem[3374] = 'd184;
    mem[3375] = 'd228;
    mem[3376] = 'd156;
    mem[3377] = 'd192;
    mem[3378] = 'd204;
    mem[3379] = 'd260;
    mem[3380] = 'd336;
    mem[3381] = 'd432;
    mem[3382] = 'd636;
    mem[3383] = 'd804;
    mem[3384] = 'd828;
    mem[3385] = 'd1004;
    mem[3386] = 'd856;
    mem[3387] = 'd1020;
    mem[3388] = 'd864;
    mem[3389] = 'd1020;
    mem[3390] = 'd864;
    mem[3391] = 'd1020;
    mem[3392] = 'd864;
    mem[3393] = 'd1020;
    mem[3394] = 'd864;
    mem[3395] = 'd1020;
    mem[3396] = 'd856;
    mem[3397] = 'd1016;
    mem[3398] = 'd812;
    mem[3399] = 'd996;
    mem[3400] = 'd572;
    mem[3401] = 'd736;
    mem[3402] = 'd292;
    mem[3403] = 'd376;
    mem[3404] = 'd188;
    mem[3405] = 'd244;
    mem[3406] = 'd148;
    mem[3407] = 'd188;
    mem[3408] = 'd176;
    mem[3409] = 'd232;
    mem[3410] = 'd276;
    mem[3411] = 'd384;
    mem[3412] = 'd428;
    mem[3413] = 'd604;
    mem[3414] = 'd632;
    mem[3415] = 'd900;
    mem[3416] = 'd692;
    mem[3417] = 'd956;
    mem[3418] = 'd724;
    mem[3419] = 'd1004;
    mem[3420] = 'd700;
    mem[3421] = 'd1004;
    mem[3422] = 'd636;
    mem[3423] = 'd964;
    mem[3424] = 'd548;
    mem[3425] = 'd912;
    mem[3426] = 'd568;
    mem[3427] = 'd872;
    mem[3428] = 'd1020;
    mem[3429] = 'd1020;
    mem[3430] = 'd1020;
    mem[3431] = 'd1020;
    mem[3432] = 'd1020;
    mem[3433] = 'd1020;
    mem[3434] = 'd448;
    mem[3435] = 'd676;
    mem[3436] = 'd20;
    mem[3437] = 'd516;
    mem[3438] = 'd44;
    mem[3439] = 'd612;
    mem[3440] = 'd68;
    mem[3441] = 'd684;
    mem[3442] = 'd120;
    mem[3443] = 'd720;
    mem[3444] = 'd172;
    mem[3445] = 'd744;
    mem[3446] = 'd188;
    mem[3447] = 'd760;
    mem[3448] = 'd180;
    mem[3449] = 'd760;
    mem[3450] = 'd172;
    mem[3451] = 'd756;
    mem[3452] = 'd160;
    mem[3453] = 'd756;
    mem[3454] = 'd164;
    mem[3455] = 'd768;
    mem[3456] = 'd176;
    mem[3457] = 'd788;
    mem[3458] = 'd196;
    mem[3459] = 'd812;
    mem[3460] = 'd204;
    mem[3461] = 'd836;
    mem[3462] = 'd208;
    mem[3463] = 'd844;
    mem[3464] = 'd212;
    mem[3465] = 'd848;
    mem[3466] = 'd208;
    mem[3467] = 'd852;
    mem[3468] = 'd208;
    mem[3469] = 'd852;
    mem[3470] = 'd208;
    mem[3471] = 'd852;
    mem[3472] = 'd208;
    mem[3473] = 'd852;
    mem[3474] = 'd208;
    mem[3475] = 'd852;
    mem[3476] = 'd208;
    mem[3477] = 'd844;
    mem[3478] = 'd200;
    mem[3479] = 'd832;
    mem[3480] = 'd184;
    mem[3481] = 'd800;
    mem[3482] = 'd160;
    mem[3483] = 'd764;
    mem[3484] = 'd148;
    mem[3485] = 'd744;
    mem[3486] = 'd148;
    mem[3487] = 'd736;
    mem[3488] = 'd160;
    mem[3489] = 'd740;
    mem[3490] = 'd172;
    mem[3491] = 'd748;
    mem[3492] = 'd188;
    mem[3493] = 'd756;
    mem[3494] = 'd172;
    mem[3495] = 'd748;
    mem[3496] = 'd120;
    mem[3497] = 'd724;
    mem[3498] = 'd72;
    mem[3499] = 'd684;
    mem[3500] = 'd48;
    mem[3501] = 'd616;
    mem[3502] = 'd24;
    mem[3503] = 'd524;
    mem[3504] = 'd404;
    mem[3505] = 'd660;
    mem[3506] = 'd1020;
    mem[3507] = 'd1020;
    mem[3508] = 'd1020;
    mem[3509] = 'd1020;
    mem[3510] = 'd1020;
    mem[3511] = 'd1020;
    mem[3512] = 'd676;
    mem[3513] = 'd900;
    mem[3514] = 'd516;
    mem[3515] = 'd884;
    mem[3516] = 'd612;
    mem[3517] = 'd944;
    mem[3518] = 'd684;
    mem[3519] = 'd996;
    mem[3520] = 'd720;
    mem[3521] = 'd1012;
    mem[3522] = 'd744;
    mem[3523] = 'd1016;
    mem[3524] = 'd760;
    mem[3525] = 'd1012;
    mem[3526] = 'd760;
    mem[3527] = 'd1000;
    mem[3528] = 'd756;
    mem[3529] = 'd988;
    mem[3530] = 'd756;
    mem[3531] = 'd988;
    mem[3532] = 'd768;
    mem[3533] = 'd992;
    mem[3534] = 'd788;
    mem[3535] = 'd1000;
    mem[3536] = 'd812;
    mem[3537] = 'd1008;
    mem[3538] = 'd836;
    mem[3539] = 'd1016;
    mem[3540] = 'd844;
    mem[3541] = 'd1020;
    mem[3542] = 'd848;
    mem[3543] = 'd1020;
    mem[3544] = 'd852;
    mem[3545] = 'd1020;
    mem[3546] = 'd852;
    mem[3547] = 'd1020;
    mem[3548] = 'd852;
    mem[3549] = 'd1020;
    mem[3550] = 'd852;
    mem[3551] = 'd1020;
    mem[3552] = 'd852;
    mem[3553] = 'd1020;
    mem[3554] = 'd844;
    mem[3555] = 'd1020;
    mem[3556] = 'd832;
    mem[3557] = 'd1012;
    mem[3558] = 'd800;
    mem[3559] = 'd996;
    mem[3560] = 'd764;
    mem[3561] = 'd984;
    mem[3562] = 'd744;
    mem[3563] = 'd976;
    mem[3564] = 'd736;
    mem[3565] = 'd972;
    mem[3566] = 'd740;
    mem[3567] = 'd976;
    mem[3568] = 'd748;
    mem[3569] = 'd992;
    mem[3570] = 'd756;
    mem[3571] = 'd1008;
    mem[3572] = 'd748;
    mem[3573] = 'd1016;
    mem[3574] = 'd724;
    mem[3575] = 'd1012;
    mem[3576] = 'd684;
    mem[3577] = 'd996;
    mem[3578] = 'd616;
    mem[3579] = 'd948;
    mem[3580] = 'd524;
    mem[3581] = 'd892;
    mem[3582] = 'd660;
    mem[3583] = 'd892;
    mem[3584] = 'd1020;
    mem[3585] = 'd1020;
    mem[3586] = 'd1020;
    mem[3587] = 'd1020;
    mem[3588] = 'd1020;
    mem[3589] = 'd1020;
    mem[3590] = 'd676;
    mem[3591] = 'd808;
    mem[3592] = 'd16;
    mem[3593] = 'd488;
    mem[3594] = 'd40;
    mem[3595] = 'd584;
    mem[3596] = 'd64;
    mem[3597] = 'd660;
    mem[3598] = 'd92;
    mem[3599] = 'd704;
    mem[3600] = 'd140;
    mem[3601] = 'd732;
    mem[3602] = 'd184;
    mem[3603] = 'd756;
    mem[3604] = 'd208;
    mem[3605] = 'd772;
    mem[3606] = 'd212;
    mem[3607] = 'd784;
    mem[3608] = 'd200;
    mem[3609] = 'd780;
    mem[3610] = 'd204;
    mem[3611] = 'd800;
    mem[3612] = 'd212;
    mem[3613] = 'd816;
    mem[3614] = 'd216;
    mem[3615] = 'd824;
    mem[3616] = 'd216;
    mem[3617] = 'd832;
    mem[3618] = 'd216;
    mem[3619] = 'd836;
    mem[3620] = 'd216;
    mem[3621] = 'd836;
    mem[3622] = 'd216;
    mem[3623] = 'd840;
    mem[3624] = 'd220;
    mem[3625] = 'd840;
    mem[3626] = 'd216;
    mem[3627] = 'd844;
    mem[3628] = 'd216;
    mem[3629] = 'd840;
    mem[3630] = 'd216;
    mem[3631] = 'd836;
    mem[3632] = 'd216;
    mem[3633] = 'd836;
    mem[3634] = 'd216;
    mem[3635] = 'd832;
    mem[3636] = 'd216;
    mem[3637] = 'd824;
    mem[3638] = 'd216;
    mem[3639] = 'd820;
    mem[3640] = 'd208;
    mem[3641] = 'd800;
    mem[3642] = 'd200;
    mem[3643] = 'd776;
    mem[3644] = 'd212;
    mem[3645] = 'd784;
    mem[3646] = 'd208;
    mem[3647] = 'd772;
    mem[3648] = 'd184;
    mem[3649] = 'd756;
    mem[3650] = 'd144;
    mem[3651] = 'd732;
    mem[3652] = 'd92;
    mem[3653] = 'd708;
    mem[3654] = 'd64;
    mem[3655] = 'd660;
    mem[3656] = 'd44;
    mem[3657] = 'd588;
    mem[3658] = 'd16;
    mem[3659] = 'd492;
    mem[3660] = 'd636;
    mem[3661] = 'd788;
    mem[3662] = 'd1020;
    mem[3663] = 'd1020;
    mem[3664] = 'd1020;
    mem[3665] = 'd1020;
    mem[3666] = 'd1020;
    mem[3667] = 'd1020;
    mem[3668] = 'd808;
    mem[3669] = 'd936;
    mem[3670] = 'd488;
    mem[3671] = 'd860;
    mem[3672] = 'd584;
    mem[3673] = 'd924;
    mem[3674] = 'd660;
    mem[3675] = 'd976;
    mem[3676] = 'd704;
    mem[3677] = 'd1008;
    mem[3678] = 'd732;
    mem[3679] = 'd1016;
    mem[3680] = 'd756;
    mem[3681] = 'd1020;
    mem[3682] = 'd772;
    mem[3683] = 'd1020;
    mem[3684] = 'd784;
    mem[3685] = 'd1020;
    mem[3686] = 'd780;
    mem[3687] = 'd1008;
    mem[3688] = 'd800;
    mem[3689] = 'd1012;
    mem[3690] = 'd816;
    mem[3691] = 'd1020;
    mem[3692] = 'd824;
    mem[3693] = 'd1020;
    mem[3694] = 'd832;
    mem[3695] = 'd1020;
    mem[3696] = 'd836;
    mem[3697] = 'd1020;
    mem[3698] = 'd836;
    mem[3699] = 'd1020;
    mem[3700] = 'd840;
    mem[3701] = 'd1020;
    mem[3702] = 'd840;
    mem[3703] = 'd1020;
    mem[3704] = 'd844;
    mem[3705] = 'd1020;
    mem[3706] = 'd840;
    mem[3707] = 'd1020;
    mem[3708] = 'd836;
    mem[3709] = 'd1020;
    mem[3710] = 'd836;
    mem[3711] = 'd1020;
    mem[3712] = 'd832;
    mem[3713] = 'd1020;
    mem[3714] = 'd824;
    mem[3715] = 'd1020;
    mem[3716] = 'd820;
    mem[3717] = 'd1020;
    mem[3718] = 'd800;
    mem[3719] = 'd1016;
    mem[3720] = 'd776;
    mem[3721] = 'd1012;
    mem[3722] = 'd784;
    mem[3723] = 'd1020;
    mem[3724] = 'd772;
    mem[3725] = 'd1020;
    mem[3726] = 'd756;
    mem[3727] = 'd1020;
    mem[3728] = 'd732;
    mem[3729] = 'd1016;
    mem[3730] = 'd708;
    mem[3731] = 'd1008;
    mem[3732] = 'd660;
    mem[3733] = 'd976;
    mem[3734] = 'd588;
    mem[3735] = 'd928;
    mem[3736] = 'd492;
    mem[3737] = 'd864;
    mem[3738] = 'd788;
    mem[3739] = 'd928;
    mem[3740] = 'd1020;
    mem[3741] = 'd1020;
    mem[3742] = 'd1020;
    mem[3743] = 'd1020;
    mem[3744] = 'd1020;
    mem[3745] = 'd1020;
    mem[3746] = 'd944;
    mem[3747] = 'd968;
    mem[3748] = 'd36;
    mem[3749] = 'd460;
    mem[3750] = 'd36;
    mem[3751] = 'd548;
    mem[3752] = 'd56;
    mem[3753] = 'd636;
    mem[3754] = 'd76;
    mem[3755] = 'd684;
    mem[3756] = 'd108;
    mem[3757] = 'd716;
    mem[3758] = 'd156;
    mem[3759] = 'd740;
    mem[3760] = 'd196;
    mem[3761] = 'd756;
    mem[3762] = 'd216;
    mem[3763] = 'd772;
    mem[3764] = 'd112;
    mem[3765] = 'd480;
    mem[3766] = 'd104;
    mem[3767] = 'd500;
    mem[3768] = 'd200;
    mem[3769] = 'd776;
    mem[3770] = 'd216;
    mem[3771] = 'd812;
    mem[3772] = 'd224;
    mem[3773] = 'd820;
    mem[3774] = 'd220;
    mem[3775] = 'd824;
    mem[3776] = 'd224;
    mem[3777] = 'd828;
    mem[3778] = 'd220;
    mem[3779] = 'd828;
    mem[3780] = 'd220;
    mem[3781] = 'd828;
    mem[3782] = 'd220;
    mem[3783] = 'd828;
    mem[3784] = 'd220;
    mem[3785] = 'd828;
    mem[3786] = 'd220;
    mem[3787] = 'd828;
    mem[3788] = 'd220;
    mem[3789] = 'd824;
    mem[3790] = 'd220;
    mem[3791] = 'd820;
    mem[3792] = 'd220;
    mem[3793] = 'd812;
    mem[3794] = 'd200;
    mem[3795] = 'd772;
    mem[3796] = 'd84;
    mem[3797] = 'd436;
    mem[3798] = 'd136;
    mem[3799] = 'd544;
    mem[3800] = 'd216;
    mem[3801] = 'd772;
    mem[3802] = 'd196;
    mem[3803] = 'd756;
    mem[3804] = 'd156;
    mem[3805] = 'd736;
    mem[3806] = 'd112;
    mem[3807] = 'd720;
    mem[3808] = 'd76;
    mem[3809] = 'd684;
    mem[3810] = 'd60;
    mem[3811] = 'd636;
    mem[3812] = 'd36;
    mem[3813] = 'd556;
    mem[3814] = 'd24;
    mem[3815] = 'd464;
    mem[3816] = 'd916;
    mem[3817] = 'd952;
    mem[3818] = 'd1020;
    mem[3819] = 'd1020;
    mem[3820] = 'd1020;
    mem[3821] = 'd1020;
    mem[3822] = 'd1020;
    mem[3823] = 'd1020;
    mem[3824] = 'd968;
    mem[3825] = 'd996;
    mem[3826] = 'd460;
    mem[3827] = 'd832;
    mem[3828] = 'd548;
    mem[3829] = 'd896;
    mem[3830] = 'd636;
    mem[3831] = 'd956;
    mem[3832] = 'd684;
    mem[3833] = 'd996;
    mem[3834] = 'd716;
    mem[3835] = 'd1012;
    mem[3836] = 'd740;
    mem[3837] = 'd1016;
    mem[3838] = 'd756;
    mem[3839] = 'd1020;
    mem[3840] = 'd772;
    mem[3841] = 'd1020;
    mem[3842] = 'd480;
    mem[3843] = 'd704;
    mem[3844] = 'd500;
    mem[3845] = 'd748;
    mem[3846] = 'd776;
    mem[3847] = 'd1000;
    mem[3848] = 'd812;
    mem[3849] = 'd1020;
    mem[3850] = 'd820;
    mem[3851] = 'd1020;
    mem[3852] = 'd824;
    mem[3853] = 'd1020;
    mem[3854] = 'd828;
    mem[3855] = 'd1020;
    mem[3856] = 'd828;
    mem[3857] = 'd1020;
    mem[3858] = 'd828;
    mem[3859] = 'd1020;
    mem[3860] = 'd828;
    mem[3861] = 'd1020;
    mem[3862] = 'd828;
    mem[3863] = 'd1020;
    mem[3864] = 'd828;
    mem[3865] = 'd1020;
    mem[3866] = 'd824;
    mem[3867] = 'd1020;
    mem[3868] = 'd820;
    mem[3869] = 'd1020;
    mem[3870] = 'd812;
    mem[3871] = 'd1020;
    mem[3872] = 'd772;
    mem[3873] = 'd1000;
    mem[3874] = 'd436;
    mem[3875] = 'd680;
    mem[3876] = 'd544;
    mem[3877] = 'd760;
    mem[3878] = 'd772;
    mem[3879] = 'd1020;
    mem[3880] = 'd756;
    mem[3881] = 'd1020;
    mem[3882] = 'd736;
    mem[3883] = 'd1016;
    mem[3884] = 'd720;
    mem[3885] = 'd1012;
    mem[3886] = 'd684;
    mem[3887] = 'd1000;
    mem[3888] = 'd636;
    mem[3889] = 'd956;
    mem[3890] = 'd556;
    mem[3891] = 'd904;
    mem[3892] = 'd464;
    mem[3893] = 'd840;
    mem[3894] = 'd952;
    mem[3895] = 'd984;
    mem[3896] = 'd1020;
    mem[3897] = 'd1020;
    mem[3898] = 'd1020;
    mem[3899] = 'd1020;
    mem[3900] = 'd1020;
    mem[3901] = 'd1020;
    mem[3902] = 'd1020;
    mem[3903] = 'd1020;
    mem[3904] = 'd356;
    mem[3905] = 'd624;
    mem[3906] = 'd24;
    mem[3907] = 'd504;
    mem[3908] = 'd52;
    mem[3909] = 'd600;
    mem[3910] = 'd68;
    mem[3911] = 'd656;
    mem[3912] = 'd84;
    mem[3913] = 'd692;
    mem[3914] = 'd112;
    mem[3915] = 'd720;
    mem[3916] = 'd160;
    mem[3917] = 'd740;
    mem[3918] = 'd192;
    mem[3919] = 'd756;
    mem[3920] = 'd224;
    mem[3921] = 'd736;
    mem[3922] = 'd44;
    mem[3923] = 'd288;
    mem[3924] = 'd44;
    mem[3925] = 'd332;
    mem[3926] = 'd128;
    mem[3927] = 'd572;
    mem[3928] = 'd204;
    mem[3929] = 'd764;
    mem[3930] = 'd224;
    mem[3931] = 'd804;
    mem[3932] = 'd228;
    mem[3933] = 'd812;
    mem[3934] = 'd228;
    mem[3935] = 'd812;
    mem[3936] = 'd228;
    mem[3937] = 'd816;
    mem[3938] = 'd228;
    mem[3939] = 'd816;
    mem[3940] = 'd228;
    mem[3941] = 'd812;
    mem[3942] = 'd224;
    mem[3943] = 'd808;
    mem[3944] = 'd220;
    mem[3945] = 'd796;
    mem[3946] = 'd192;
    mem[3947] = 'd736;
    mem[3948] = 'd116;
    mem[3949] = 'd532;
    mem[3950] = 'd36;
    mem[3951] = 'd300;
    mem[3952] = 'd64;
    mem[3953] = 'd328;
    mem[3954] = 'd236;
    mem[3955] = 'd772;
    mem[3956] = 'd196;
    mem[3957] = 'd752;
    mem[3958] = 'd160;
    mem[3959] = 'd740;
    mem[3960] = 'd116;
    mem[3961] = 'd724;
    mem[3962] = 'd84;
    mem[3963] = 'd696;
    mem[3964] = 'd72;
    mem[3965] = 'd660;
    mem[3966] = 'd56;
    mem[3967] = 'd604;
    mem[3968] = 'd28;
    mem[3969] = 'd508;
    mem[3970] = 'd292;
    mem[3971] = 'd584;
    mem[3972] = 'd1020;
    mem[3973] = 'd1020;
    mem[3974] = 'd1020;
    mem[3975] = 'd1020;
    mem[3976] = 'd1020;
    mem[3977] = 'd1020;
    mem[3978] = 'd1020;
    mem[3979] = 'd1020;
    mem[3980] = 'd1020;
    mem[3981] = 'd1020;
    mem[3982] = 'd624;
    mem[3983] = 'd876;
    mem[3984] = 'd504;
    mem[3985] = 'd860;
    mem[3986] = 'd600;
    mem[3987] = 'd924;
    mem[3988] = 'd656;
    mem[3989] = 'd972;
    mem[3990] = 'd692;
    mem[3991] = 'd1004;
    mem[3992] = 'd720;
    mem[3993] = 'd1016;
    mem[3994] = 'd740;
    mem[3995] = 'd1016;
    mem[3996] = 'd756;
    mem[3997] = 'd1020;
    mem[3998] = 'd736;
    mem[3999] = 'd948;
    mem[4000] = 'd288;
    mem[4001] = 'd500;
    mem[4002] = 'd332;
    mem[4003] = 'd564;
    mem[4004] = 'd572;
    mem[4005] = 'd820;
    mem[4006] = 'd764;
    mem[4007] = 'd1000;
    mem[4008] = 'd804;
    mem[4009] = 'd1016;
    mem[4010] = 'd812;
    mem[4011] = 'd1020;
    mem[4012] = 'd812;
    mem[4013] = 'd1020;
    mem[4014] = 'd816;
    mem[4015] = 'd1020;
    mem[4016] = 'd816;
    mem[4017] = 'd1020;
    mem[4018] = 'd812;
    mem[4019] = 'd1020;
    mem[4020] = 'd808;
    mem[4021] = 'd1020;
    mem[4022] = 'd796;
    mem[4023] = 'd1016;
    mem[4024] = 'd736;
    mem[4025] = 'd972;
    mem[4026] = 'd532;
    mem[4027] = 'd780;
    mem[4028] = 'd300;
    mem[4029] = 'd528;
    mem[4030] = 'd328;
    mem[4031] = 'd528;
    mem[4032] = 'd772;
    mem[4033] = 'd988;
    mem[4034] = 'd752;
    mem[4035] = 'd1020;
    mem[4036] = 'd740;
    mem[4037] = 'd1016;
    mem[4038] = 'd724;
    mem[4039] = 'd1016;
    mem[4040] = 'd696;
    mem[4041] = 'd1004;
    mem[4042] = 'd660;
    mem[4043] = 'd972;
    mem[4044] = 'd604;
    mem[4045] = 'd928;
    mem[4046] = 'd508;
    mem[4047] = 'd868;
    mem[4048] = 'd584;
    mem[4049] = 'd864;
    mem[4050] = 'd1020;
    mem[4051] = 'd1020;
    mem[4052] = 'd1020;
    mem[4053] = 'd1020;
    mem[4054] = 'd1020;
    mem[4055] = 'd1020;
    mem[4056] = 'd1020;
    mem[4057] = 'd1020;
    mem[4058] = 'd1020;
    mem[4059] = 'd1020;
    mem[4060] = 'd792;
    mem[4061] = 'd876;
    mem[4062] = 'd12;
    mem[4063] = 'd456;
    mem[4064] = 'd40;
    mem[4065] = 'd556;
    mem[4066] = 'd64;
    mem[4067] = 'd624;
    mem[4068] = 'd80;
    mem[4069] = 'd668;
    mem[4070] = 'd88;
    mem[4071] = 'd700;
    mem[4072] = 'd116;
    mem[4073] = 'd716;
    mem[4074] = 'd156;
    mem[4075] = 'd736;
    mem[4076] = 'd192;
    mem[4077] = 'd752;
    mem[4078] = 'd216;
    mem[4079] = 'd712;
    mem[4080] = 'd48;
    mem[4081] = 'd332;
    mem[4082] = 'd20;
    mem[4083] = 'd252;
    mem[4084] = 'd32;
    mem[4085] = 'd288;
    mem[4086] = 'd76;
    mem[4087] = 'd420;
    mem[4088] = 'd120;
    mem[4089] = 'd548;
    mem[4090] = 'd152;
    mem[4091] = 'd640;
    mem[4092] = 'd168;
    mem[4093] = 'd676;
    mem[4094] = 'd164;
    mem[4095] = 'd672;
    mem[4096] = 'd152;
    mem[4097] = 'd628;
    mem[4098] = 'd116;
    mem[4099] = 'd536;
    mem[4100] = 'd72;
    mem[4101] = 'd404;
    mem[4102] = 'd32;
    mem[4103] = 'd288;
    mem[4104] = 'd16;
    mem[4105] = 'd256;
    mem[4106] = 'd68;
    mem[4107] = 'd372;
    mem[4108] = 'd232;
    mem[4109] = 'd752;
    mem[4110] = 'd188;
    mem[4111] = 'd752;
    mem[4112] = 'd156;
    mem[4113] = 'd736;
    mem[4114] = 'd116;
    mem[4115] = 'd720;
    mem[4116] = 'd92;
    mem[4117] = 'd696;
    mem[4118] = 'd80;
    mem[4119] = 'd668;
    mem[4120] = 'd68;
    mem[4121] = 'd628;
    mem[4122] = 'd44;
    mem[4123] = 'd556;
    mem[4124] = 'd20;
    mem[4125] = 'd464;
    mem[4126] = 'd744;
    mem[4127] = 'd848;
    mem[4128] = 'd1020;
    mem[4129] = 'd1020;
    mem[4130] = 'd1020;
    mem[4131] = 'd1020;
    mem[4132] = 'd1020;
    mem[4133] = 'd1020;
    mem[4134] = 'd1020;
    mem[4135] = 'd1020;
    mem[4136] = 'd1020;
    mem[4137] = 'd1020;
    mem[4138] = 'd876;
    mem[4139] = 'd956;
    mem[4140] = 'd456;
    mem[4141] = 'd836;
    mem[4142] = 'd556;
    mem[4143] = 'd892;
    mem[4144] = 'd624;
    mem[4145] = 'd940;
    mem[4146] = 'd668;
    mem[4147] = 'd980;
    mem[4148] = 'd700;
    mem[4149] = 'd1008;
    mem[4150] = 'd716;
    mem[4151] = 'd1016;
    mem[4152] = 'd736;
    mem[4153] = 'd1020;
    mem[4154] = 'd752;
    mem[4155] = 'd1020;
    mem[4156] = 'd712;
    mem[4157] = 'd912;
    mem[4158] = 'd332;
    mem[4159] = 'd552;
    mem[4160] = 'd252;
    mem[4161] = 'd476;
    mem[4162] = 'd288;
    mem[4163] = 'd520;
    mem[4164] = 'd420;
    mem[4165] = 'd668;
    mem[4166] = 'd548;
    mem[4167] = 'd804;
    mem[4168] = 'd640;
    mem[4169] = 'd892;
    mem[4170] = 'd676;
    mem[4171] = 'd928;
    mem[4172] = 'd672;
    mem[4173] = 'd924;
    mem[4174] = 'd628;
    mem[4175] = 'd880;
    mem[4176] = 'd536;
    mem[4177] = 'd788;
    mem[4178] = 'd404;
    mem[4179] = 'd652;
    mem[4180] = 'd288;
    mem[4181] = 'd516;
    mem[4182] = 'd256;
    mem[4183] = 'd480;
    mem[4184] = 'd372;
    mem[4185] = 'd584;
    mem[4186] = 'd752;
    mem[4187] = 'd956;
    mem[4188] = 'd752;
    mem[4189] = 'd1020;
    mem[4190] = 'd736;
    mem[4191] = 'd1020;
    mem[4192] = 'd720;
    mem[4193] = 'd1016;
    mem[4194] = 'd696;
    mem[4195] = 'd1008;
    mem[4196] = 'd668;
    mem[4197] = 'd980;
    mem[4198] = 'd628;
    mem[4199] = 'd948;
    mem[4200] = 'd556;
    mem[4201] = 'd892;
    mem[4202] = 'd464;
    mem[4203] = 'd836;
    mem[4204] = 'd848;
    mem[4205] = 'd952;
    mem[4206] = 'd1020;
    mem[4207] = 'd1020;
    mem[4208] = 'd1020;
    mem[4209] = 'd1020;
    mem[4210] = 'd1020;
    mem[4211] = 'd1020;
    mem[4212] = 'd1020;
    mem[4213] = 'd1020;
    mem[4214] = 'd1020;
    mem[4215] = 'd1020;
    mem[4216] = 'd1020;
    mem[4217] = 'd1020;
    mem[4218] = 'd280;
    mem[4219] = 'd576;
    mem[4220] = 'd28;
    mem[4221] = 'd504;
    mem[4222] = 'd52;
    mem[4223] = 'd580;
    mem[4224] = 'd72;
    mem[4225] = 'd636;
    mem[4226] = 'd84;
    mem[4227] = 'd672;
    mem[4228] = 'd92;
    mem[4229] = 'd696;
    mem[4230] = 'd108;
    mem[4231] = 'd716;
    mem[4232] = 'd144;
    mem[4233] = 'd732;
    mem[4234] = 'd180;
    mem[4235] = 'd748;
    mem[4236] = 'd224;
    mem[4237] = 'd752;
    mem[4238] = 'd112;
    mem[4239] = 'd480;
    mem[4240] = 'd20;
    mem[4241] = 'd308;
    mem[4242] = 'd20;
    mem[4243] = 'd296;
    mem[4244] = 'd16;
    mem[4245] = 'd264;
    mem[4246] = 'd20;
    mem[4247] = 'd248;
    mem[4248] = 'd20;
    mem[4249] = 'd244;
    mem[4250] = 'd20;
    mem[4251] = 'd248;
    mem[4252] = 'd20;
    mem[4253] = 'd252;
    mem[4254] = 'd16;
    mem[4255] = 'd268;
    mem[4256] = 'd20;
    mem[4257] = 'd300;
    mem[4258] = 'd28;
    mem[4259] = 'd328;
    mem[4260] = 'd136;
    mem[4261] = 'd532;
    mem[4262] = 'd224;
    mem[4263] = 'd768;
    mem[4264] = 'd176;
    mem[4265] = 'd748;
    mem[4266] = 'd144;
    mem[4267] = 'd732;
    mem[4268] = 'd112;
    mem[4269] = 'd716;
    mem[4270] = 'd92;
    mem[4271] = 'd696;
    mem[4272] = 'd84;
    mem[4273] = 'd676;
    mem[4274] = 'd76;
    mem[4275] = 'd640;
    mem[4276] = 'd56;
    mem[4277] = 'd588;
    mem[4278] = 'd32;
    mem[4279] = 'd508;
    mem[4280] = 'd256;
    mem[4281] = 'd564;
    mem[4282] = 'd1008;
    mem[4283] = 'd1012;
    mem[4284] = 'd1020;
    mem[4285] = 'd1020;
    mem[4286] = 'd1020;
    mem[4287] = 'd1020;
    mem[4288] = 'd1020;
    mem[4289] = 'd1020;
    mem[4290] = 'd1020;
    mem[4291] = 'd1020;
    mem[4292] = 'd1020;
    mem[4293] = 'd1020;
    mem[4294] = 'd1020;
    mem[4295] = 'd1020;
    mem[4296] = 'd576;
    mem[4297] = 'd856;
    mem[4298] = 'd504;
    mem[4299] = 'd856;
    mem[4300] = 'd580;
    mem[4301] = 'd904;
    mem[4302] = 'd636;
    mem[4303] = 'd952;
    mem[4304] = 'd672;
    mem[4305] = 'd984;
    mem[4306] = 'd696;
    mem[4307] = 'd1004;
    mem[4308] = 'd716;
    mem[4309] = 'd1020;
    mem[4310] = 'd732;
    mem[4311] = 'd1020;
    mem[4312] = 'd748;
    mem[4313] = 'd1020;
    mem[4314] = 'd752;
    mem[4315] = 'd956;
    mem[4316] = 'd480;
    mem[4317] = 'd680;
    mem[4318] = 'd308;
    mem[4319] = 'd544;
    mem[4320] = 'd296;
    mem[4321] = 'd528;
    mem[4322] = 'd264;
    mem[4323] = 'd488;
    mem[4324] = 'd248;
    mem[4325] = 'd468;
    mem[4326] = 'd244;
    mem[4327] = 'd468;
    mem[4328] = 'd248;
    mem[4329] = 'd468;
    mem[4330] = 'd252;
    mem[4331] = 'd472;
    mem[4332] = 'd268;
    mem[4333] = 'd496;
    mem[4334] = 'd300;
    mem[4335] = 'd528;
    mem[4336] = 'd328;
    mem[4337] = 'd560;
    mem[4338] = 'd532;
    mem[4339] = 'd728;
    mem[4340] = 'd768;
    mem[4341] = 'd976;
    mem[4342] = 'd748;
    mem[4343] = 'd1020;
    mem[4344] = 'd732;
    mem[4345] = 'd1020;
    mem[4346] = 'd716;
    mem[4347] = 'd1020;
    mem[4348] = 'd696;
    mem[4349] = 'd1008;
    mem[4350] = 'd676;
    mem[4351] = 'd984;
    mem[4352] = 'd640;
    mem[4353] = 'd956;
    mem[4354] = 'd588;
    mem[4355] = 'd912;
    mem[4356] = 'd508;
    mem[4357] = 'd860;
    mem[4358] = 'd564;
    mem[4359] = 'd856;
    mem[4360] = 'd1012;
    mem[4361] = 'd1012;
    mem[4362] = 'd1020;
    mem[4363] = 'd1020;
    mem[4364] = 'd1020;
    mem[4365] = 'd1020;
    mem[4366] = 'd1020;
    mem[4367] = 'd1020;
    mem[4368] = 'd1020;
    mem[4369] = 'd1020;
    mem[4370] = 'd1020;
    mem[4371] = 'd1020;
    mem[4372] = 'd1020;
    mem[4373] = 'd1020;
    mem[4374] = 'd848;
    mem[4375] = 'd912;
    mem[4376] = 'd24;
    mem[4377] = 'd456;
    mem[4378] = 'd36;
    mem[4379] = 'd528;
    mem[4380] = 'd60;
    mem[4381] = 'd596;
    mem[4382] = 'd76;
    mem[4383] = 'd640;
    mem[4384] = 'd88;
    mem[4385] = 'd672;
    mem[4386] = 'd92;
    mem[4387] = 'd692;
    mem[4388] = 'd100;
    mem[4389] = 'd708;
    mem[4390] = 'd124;
    mem[4391] = 'd724;
    mem[4392] = 'd152;
    mem[4393] = 'd736;
    mem[4394] = 'd200;
    mem[4395] = 'd768;
    mem[4396] = 'd204;
    mem[4397] = 'd708;
    mem[4398] = 'd132;
    mem[4399] = 'd532;
    mem[4400] = 'd60;
    mem[4401] = 'd400;
    mem[4402] = 'd32;
    mem[4403] = 'd352;
    mem[4404] = 'd24;
    mem[4405] = 'd344;
    mem[4406] = 'd28;
    mem[4407] = 'd344;
    mem[4408] = 'd36;
    mem[4409] = 'd364;
    mem[4410] = 'd72;
    mem[4411] = 'd420;
    mem[4412] = 'd140;
    mem[4413] = 'd556;
    mem[4414] = 'd204;
    mem[4415] = 'd716;
    mem[4416] = 'd192;
    mem[4417] = 'd764;
    mem[4418] = 'd156;
    mem[4419] = 'd736;
    mem[4420] = 'd128;
    mem[4421] = 'd724;
    mem[4422] = 'd100;
    mem[4423] = 'd708;
    mem[4424] = 'd92;
    mem[4425] = 'd692;
    mem[4426] = 'd88;
    mem[4427] = 'd672;
    mem[4428] = 'd80;
    mem[4429] = 'd644;
    mem[4430] = 'd64;
    mem[4431] = 'd600;
    mem[4432] = 'd40;
    mem[4433] = 'd532;
    mem[4434] = 'd52;
    mem[4435] = 'd472;
    mem[4436] = 'd796;
    mem[4437] = 'd880;
    mem[4438] = 'd1020;
    mem[4439] = 'd1020;
    mem[4440] = 'd1020;
    mem[4441] = 'd1020;
    mem[4442] = 'd1020;
    mem[4443] = 'd1020;
    mem[4444] = 'd1020;
    mem[4445] = 'd1020;
    mem[4446] = 'd1020;
    mem[4447] = 'd1020;
    mem[4448] = 'd1020;
    mem[4449] = 'd1020;
    mem[4450] = 'd1020;
    mem[4451] = 'd1020;
    mem[4452] = 'd912;
    mem[4453] = 'd972;
    mem[4454] = 'd456;
    mem[4455] = 'd828;
    mem[4456] = 'd528;
    mem[4457] = 'd868;
    mem[4458] = 'd596;
    mem[4459] = 'd916;
    mem[4460] = 'd640;
    mem[4461] = 'd956;
    mem[4462] = 'd672;
    mem[4463] = 'd984;
    mem[4464] = 'd692;
    mem[4465] = 'd1004;
    mem[4466] = 'd708;
    mem[4467] = 'd1016;
    mem[4468] = 'd724;
    mem[4469] = 'd1020;
    mem[4470] = 'd736;
    mem[4471] = 'd1020;
    mem[4472] = 'd768;
    mem[4473] = 'd1016;
    mem[4474] = 'd708;
    mem[4475] = 'd896;
    mem[4476] = 'd532;
    mem[4477] = 'd728;
    mem[4478] = 'd400;
    mem[4479] = 'd624;
    mem[4480] = 'd352;
    mem[4481] = 'd584;
    mem[4482] = 'd344;
    mem[4483] = 'd576;
    mem[4484] = 'd344;
    mem[4485] = 'd580;
    mem[4486] = 'd364;
    mem[4487] = 'd596;
    mem[4488] = 'd420;
    mem[4489] = 'd640;
    mem[4490] = 'd556;
    mem[4491] = 'd752;
    mem[4492] = 'd716;
    mem[4493] = 'd916;
    mem[4494] = 'd764;
    mem[4495] = 'd1020;
    mem[4496] = 'd736;
    mem[4497] = 'd1020;
    mem[4498] = 'd724;
    mem[4499] = 'd1020;
    mem[4500] = 'd708;
    mem[4501] = 'd1016;
    mem[4502] = 'd692;
    mem[4503] = 'd1008;
    mem[4504] = 'd672;
    mem[4505] = 'd988;
    mem[4506] = 'd644;
    mem[4507] = 'd956;
    mem[4508] = 'd600;
    mem[4509] = 'd920;
    mem[4510] = 'd532;
    mem[4511] = 'd872;
    mem[4512] = 'd472;
    mem[4513] = 'd836;
    mem[4514] = 'd880;
    mem[4515] = 'd964;
    mem[4516] = 'd1020;
    mem[4517] = 'd1020;
    mem[4518] = 'd1020;
    mem[4519] = 'd1020;
    mem[4520] = 'd1020;
    mem[4521] = 'd1020;
    mem[4522] = 'd1020;
    mem[4523] = 'd1020;
    mem[4524] = 'd1020;
    mem[4525] = 'd1020;
    mem[4526] = 'd1020;
    mem[4527] = 'd1020;
    mem[4528] = 'd1020;
    mem[4529] = 'd1020;
    mem[4530] = 'd1016;
    mem[4531] = 'd1020;
    mem[4532] = 'd424;
    mem[4533] = 'd668;
    mem[4534] = 'd20;
    mem[4535] = 'd476;
    mem[4536] = 'd40;
    mem[4537] = 'd540;
    mem[4538] = 'd60;
    mem[4539] = 'd600;
    mem[4540] = 'd80;
    mem[4541] = 'd640;
    mem[4542] = 'd88;
    mem[4543] = 'd664;
    mem[4544] = 'd92;
    mem[4545] = 'd684;
    mem[4546] = 'd96;
    mem[4547] = 'd700;
    mem[4548] = 'd108;
    mem[4549] = 'd712;
    mem[4550] = 'd124;
    mem[4551] = 'd720;
    mem[4552] = 'd144;
    mem[4553] = 'd732;
    mem[4554] = 'd176;
    mem[4555] = 'd752;
    mem[4556] = 'd208;
    mem[4557] = 'd780;
    mem[4558] = 'd216;
    mem[4559] = 'd776;
    mem[4560] = 'd212;
    mem[4561] = 'd756;
    mem[4562] = 'd216;
    mem[4563] = 'd756;
    mem[4564] = 'd212;
    mem[4565] = 'd768;
    mem[4566] = 'd204;
    mem[4567] = 'd776;
    mem[4568] = 'd172;
    mem[4569] = 'd752;
    mem[4570] = 'd144;
    mem[4571] = 'd732;
    mem[4572] = 'd124;
    mem[4573] = 'd720;
    mem[4574] = 'd112;
    mem[4575] = 'd712;
    mem[4576] = 'd100;
    mem[4577] = 'd700;
    mem[4578] = 'd92;
    mem[4579] = 'd684;
    mem[4580] = 'd88;
    mem[4581] = 'd668;
    mem[4582] = 'd80;
    mem[4583] = 'd640;
    mem[4584] = 'd64;
    mem[4585] = 'd604;
    mem[4586] = 'd44;
    mem[4587] = 'd548;
    mem[4588] = 'd20;
    mem[4589] = 'd480;
    mem[4590] = 'd408;
    mem[4591] = 'd660;
    mem[4592] = 'd1016;
    mem[4593] = 'd1020;
    mem[4594] = 'd1020;
    mem[4595] = 'd1020;
    mem[4596] = 'd1020;
    mem[4597] = 'd1020;
    mem[4598] = 'd1020;
    mem[4599] = 'd1020;
    mem[4600] = 'd1020;
    mem[4601] = 'd1020;
    mem[4602] = 'd1020;
    mem[4603] = 'd1020;
    mem[4604] = 'd1020;
    mem[4605] = 'd1020;
    mem[4606] = 'd1020;
    mem[4607] = 'd1020;
    mem[4608] = 'd1020;
    mem[4609] = 'd1020;
    mem[4610] = 'd668;
    mem[4611] = 'd896;
    mem[4612] = 'd476;
    mem[4613] = 'd844;
    mem[4614] = 'd540;
    mem[4615] = 'd876;
    mem[4616] = 'd600;
    mem[4617] = 'd920;
    mem[4618] = 'd640;
    mem[4619] = 'd956;
    mem[4620] = 'd664;
    mem[4621] = 'd980;
    mem[4622] = 'd684;
    mem[4623] = 'd996;
    mem[4624] = 'd700;
    mem[4625] = 'd1012;
    mem[4626] = 'd712;
    mem[4627] = 'd1020;
    mem[4628] = 'd720;
    mem[4629] = 'd1020;
    mem[4630] = 'd732;
    mem[4631] = 'd1020;
    mem[4632] = 'd752;
    mem[4633] = 'd1020;
    mem[4634] = 'd780;
    mem[4635] = 'd1012;
    mem[4636] = 'd776;
    mem[4637] = 'd984;
    mem[4638] = 'd756;
    mem[4639] = 'd960;
    mem[4640] = 'd756;
    mem[4641] = 'd960;
    mem[4642] = 'd768;
    mem[4643] = 'd976;
    mem[4644] = 'd776;
    mem[4645] = 'd1012;
    mem[4646] = 'd752;
    mem[4647] = 'd1020;
    mem[4648] = 'd732;
    mem[4649] = 'd1020;
    mem[4650] = 'd720;
    mem[4651] = 'd1020;
    mem[4652] = 'd712;
    mem[4653] = 'd1020;
    mem[4654] = 'd700;
    mem[4655] = 'd1012;
    mem[4656] = 'd684;
    mem[4657] = 'd1000;
    mem[4658] = 'd668;
    mem[4659] = 'd984;
    mem[4660] = 'd640;
    mem[4661] = 'd956;
    mem[4662] = 'd604;
    mem[4663] = 'd924;
    mem[4664] = 'd548;
    mem[4665] = 'd880;
    mem[4666] = 'd480;
    mem[4667] = 'd844;
    mem[4668] = 'd660;
    mem[4669] = 'd892;
    mem[4670] = 'd1020;
    mem[4671] = 'd1020;
    mem[4672] = 'd1020;
    mem[4673] = 'd1020;
    mem[4674] = 'd1020;
    mem[4675] = 'd1020;
    mem[4676] = 'd1020;
    mem[4677] = 'd1020;
    mem[4678] = 'd1020;
    mem[4679] = 'd1020;
    mem[4680] = 'd1020;
    mem[4681] = 'd1020;
    mem[4682] = 'd1020;
    mem[4683] = 'd1020;
    mem[4684] = 'd1020;
    mem[4685] = 'd1020;
    mem[4686] = 'd1016;
    mem[4687] = 'd1020;
    mem[4688] = 'd948;
    mem[4689] = 'd976;
    mem[4690] = 'd220;
    mem[4691] = 'd540;
    mem[4692] = 'd24;
    mem[4693] = 'd488;
    mem[4694] = 'd44;
    mem[4695] = 'd548;
    mem[4696] = 'd60;
    mem[4697] = 'd596;
    mem[4698] = 'd76;
    mem[4699] = 'd632;
    mem[4700] = 'd84;
    mem[4701] = 'd656;
    mem[4702] = 'd88;
    mem[4703] = 'd672;
    mem[4704] = 'd92;
    mem[4705] = 'd688;
    mem[4706] = 'd96;
    mem[4707] = 'd696;
    mem[4708] = 'd104;
    mem[4709] = 'd704;
    mem[4710] = 'd116;
    mem[4711] = 'd712;
    mem[4712] = 'd128;
    mem[4713] = 'd716;
    mem[4714] = 'd132;
    mem[4715] = 'd716;
    mem[4716] = 'd132;
    mem[4717] = 'd720;
    mem[4718] = 'd132;
    mem[4719] = 'd716;
    mem[4720] = 'd132;
    mem[4721] = 'd716;
    mem[4722] = 'd128;
    mem[4723] = 'd716;
    mem[4724] = 'd120;
    mem[4725] = 'd712;
    mem[4726] = 'd104;
    mem[4727] = 'd704;
    mem[4728] = 'd92;
    mem[4729] = 'd696;
    mem[4730] = 'd92;
    mem[4731] = 'd688;
    mem[4732] = 'd88;
    mem[4733] = 'd676;
    mem[4734] = 'd88;
    mem[4735] = 'd660;
    mem[4736] = 'd80;
    mem[4737] = 'd636;
    mem[4738] = 'd68;
    mem[4739] = 'd600;
    mem[4740] = 'd48;
    mem[4741] = 'd552;
    mem[4742] = 'd24;
    mem[4743] = 'd492;
    mem[4744] = 'd192;
    mem[4745] = 'd520;
    mem[4746] = 'd936;
    mem[4747] = 'd964;
    mem[4748] = 'd1016;
    mem[4749] = 'd1020;
    mem[4750] = 'd1020;
    mem[4751] = 'd1020;
    mem[4752] = 'd1020;
    mem[4753] = 'd1020;
    mem[4754] = 'd1020;
    mem[4755] = 'd1020;
    mem[4756] = 'd1020;
    mem[4757] = 'd1020;
    mem[4758] = 'd1020;
    mem[4759] = 'd1020;
    mem[4760] = 'd1020;
    mem[4761] = 'd1020;
    mem[4762] = 'd1020;
    mem[4763] = 'd1020;
    mem[4764] = 'd1020;
    mem[4765] = 'd1020;
    mem[4766] = 'd976;
    mem[4767] = 'd1000;
    mem[4768] = 'd540;
    mem[4769] = 'd844;
    mem[4770] = 'd488;
    mem[4771] = 'd848;
    mem[4772] = 'd548;
    mem[4773] = 'd880;
    mem[4774] = 'd596;
    mem[4775] = 'd916;
    mem[4776] = 'd632;
    mem[4777] = 'd952;
    mem[4778] = 'd656;
    mem[4779] = 'd972;
    mem[4780] = 'd672;
    mem[4781] = 'd992;
    mem[4782] = 'd688;
    mem[4783] = 'd1004;
    mem[4784] = 'd696;
    mem[4785] = 'd1016;
    mem[4786] = 'd704;
    mem[4787] = 'd1020;
    mem[4788] = 'd712;
    mem[4789] = 'd1020;
    mem[4790] = 'd716;
    mem[4791] = 'd1020;
    mem[4792] = 'd716;
    mem[4793] = 'd1020;
    mem[4794] = 'd720;
    mem[4795] = 'd1020;
    mem[4796] = 'd716;
    mem[4797] = 'd1020;
    mem[4798] = 'd716;
    mem[4799] = 'd1020;
    mem[4800] = 'd716;
    mem[4801] = 'd1020;
    mem[4802] = 'd712;
    mem[4803] = 'd1020;
    mem[4804] = 'd704;
    mem[4805] = 'd1020;
    mem[4806] = 'd696;
    mem[4807] = 'd1016;
    mem[4808] = 'd688;
    mem[4809] = 'd1008;
    mem[4810] = 'd676;
    mem[4811] = 'd992;
    mem[4812] = 'd660;
    mem[4813] = 'd976;
    mem[4814] = 'd636;
    mem[4815] = 'd952;
    mem[4816] = 'd600;
    mem[4817] = 'd920;
    mem[4818] = 'd552;
    mem[4819] = 'd884;
    mem[4820] = 'd492;
    mem[4821] = 'd852;
    mem[4822] = 'd520;
    mem[4823] = 'd836;
    mem[4824] = 'd964;
    mem[4825] = 'd996;
    mem[4826] = 'd1020;
    mem[4827] = 'd1020;
    mem[4828] = 'd1020;
    mem[4829] = 'd1020;
    mem[4830] = 'd1020;
    mem[4831] = 'd1020;
    mem[4832] = 'd1020;
    mem[4833] = 'd1020;
    mem[4834] = 'd1020;
    mem[4835] = 'd1020;
    mem[4836] = 'd1020;
    mem[4837] = 'd1020;
    mem[4838] = 'd1020;
    mem[4839] = 'd1020;
    mem[4840] = 'd1020;
    mem[4841] = 'd1020;
    mem[4842] = 'd1020;
    mem[4843] = 'd1020;
    mem[4844] = 'd1016;
    mem[4845] = 'd1020;
    mem[4846] = 'd900;
    mem[4847] = 'd944;
    mem[4848] = 'd168;
    mem[4849] = 'd504;
    mem[4850] = 'd24;
    mem[4851] = 'd488;
    mem[4852] = 'd40;
    mem[4853] = 'd540;
    mem[4854] = 'd56;
    mem[4855] = 'd584;
    mem[4856] = 'd72;
    mem[4857] = 'd620;
    mem[4858] = 'd80;
    mem[4859] = 'd644;
    mem[4860] = 'd88;
    mem[4861] = 'd660;
    mem[4862] = 'd88;
    mem[4863] = 'd672;
    mem[4864] = 'd92;
    mem[4865] = 'd680;
    mem[4866] = 'd92;
    mem[4867] = 'd688;
    mem[4868] = 'd92;
    mem[4869] = 'd692;
    mem[4870] = 'd96;
    mem[4871] = 'd692;
    mem[4872] = 'd96;
    mem[4873] = 'd692;
    mem[4874] = 'd100;
    mem[4875] = 'd696;
    mem[4876] = 'd96;
    mem[4877] = 'd692;
    mem[4878] = 'd92;
    mem[4879] = 'd692;
    mem[4880] = 'd92;
    mem[4881] = 'd684;
    mem[4882] = 'd92;
    mem[4883] = 'd680;
    mem[4884] = 'd88;
    mem[4885] = 'd676;
    mem[4886] = 'd88;
    mem[4887] = 'd664;
    mem[4888] = 'd84;
    mem[4889] = 'd648;
    mem[4890] = 'd76;
    mem[4891] = 'd624;
    mem[4892] = 'd60;
    mem[4893] = 'd588;
    mem[4894] = 'd44;
    mem[4895] = 'd548;
    mem[4896] = 'd24;
    mem[4897] = 'd492;
    mem[4898] = 'd144;
    mem[4899] = 'd496;
    mem[4900] = 'd892;
    mem[4901] = 'd940;
    mem[4902] = 'd1016;
    mem[4903] = 'd1020;
    mem[4904] = 'd1020;
    mem[4905] = 'd1020;
    mem[4906] = 'd1020;
    mem[4907] = 'd1020;
    mem[4908] = 'd1020;
    mem[4909] = 'd1020;
    mem[4910] = 'd1020;
    mem[4911] = 'd1020;
    mem[4912] = 'd1020;
    mem[4913] = 'd1020;
    mem[4914] = 'd1020;
    mem[4915] = 'd1020;
    mem[4916] = 'd1020;
    mem[4917] = 'd1020;
    mem[4918] = 'd1020;
    mem[4919] = 'd1020;
    mem[4920] = 'd1020;
    mem[4921] = 'd1020;
    mem[4922] = 'd1020;
    mem[4923] = 'd1020;
    mem[4924] = 'd944;
    mem[4925] = 'd988;
    mem[4926] = 'd504;
    mem[4927] = 'd824;
    mem[4928] = 'd488;
    mem[4929] = 'd852;
    mem[4930] = 'd540;
    mem[4931] = 'd880;
    mem[4932] = 'd584;
    mem[4933] = 'd908;
    mem[4934] = 'd620;
    mem[4935] = 'd940;
    mem[4936] = 'd644;
    mem[4937] = 'd960;
    mem[4938] = 'd660;
    mem[4939] = 'd980;
    mem[4940] = 'd672;
    mem[4941] = 'd996;
    mem[4942] = 'd680;
    mem[4943] = 'd1004;
    mem[4944] = 'd688;
    mem[4945] = 'd1012;
    mem[4946] = 'd692;
    mem[4947] = 'd1016;
    mem[4948] = 'd692;
    mem[4949] = 'd1016;
    mem[4950] = 'd692;
    mem[4951] = 'd1016;
    mem[4952] = 'd696;
    mem[4953] = 'd1016;
    mem[4954] = 'd692;
    mem[4955] = 'd1016;
    mem[4956] = 'd692;
    mem[4957] = 'd1016;
    mem[4958] = 'd684;
    mem[4959] = 'd1012;
    mem[4960] = 'd680;
    mem[4961] = 'd1004;
    mem[4962] = 'd676;
    mem[4963] = 'd996;
    mem[4964] = 'd664;
    mem[4965] = 'd984;
    mem[4966] = 'd648;
    mem[4967] = 'd968;
    mem[4968] = 'd624;
    mem[4969] = 'd940;
    mem[4970] = 'd588;
    mem[4971] = 'd912;
    mem[4972] = 'd548;
    mem[4973] = 'd884;
    mem[4974] = 'd492;
    mem[4975] = 'd852;
    mem[4976] = 'd496;
    mem[4977] = 'd828;
    mem[4978] = 'd940;
    mem[4979] = 'd988;
    mem[4980] = 'd1020;
    mem[4981] = 'd1020;
    mem[4982] = 'd1020;
    mem[4983] = 'd1020;
    mem[4984] = 'd1020;
    mem[4985] = 'd1020;
    mem[4986] = 'd1020;
    mem[4987] = 'd1020;
    mem[4988] = 'd1020;
    mem[4989] = 'd1020;
    mem[4990] = 'd1020;
    mem[4991] = 'd1020;
    mem[4992] = 'd1020;
    mem[4993] = 'd1020;
    mem[4994] = 'd1020;
    mem[4995] = 'd1020;
    mem[4996] = 'd1020;
    mem[4997] = 'd1020;
    mem[4998] = 'd1020;
    mem[4999] = 'd1020;
    mem[5000] = 'd1016;
    mem[5001] = 'd1020;
    mem[5002] = 'd1012;
    mem[5003] = 'd1020;
    mem[5004] = 'd896;
    mem[5005] = 'd940;
    mem[5006] = 'd220;
    mem[5007] = 'd540;
    mem[5008] = 'd20;
    mem[5009] = 'd476;
    mem[5010] = 'd36;
    mem[5011] = 'd528;
    mem[5012] = 'd52;
    mem[5013] = 'd572;
    mem[5014] = 'd64;
    mem[5015] = 'd600;
    mem[5016] = 'd72;
    mem[5017] = 'd624;
    mem[5018] = 'd80;
    mem[5019] = 'd640;
    mem[5020] = 'd84;
    mem[5021] = 'd656;
    mem[5022] = 'd88;
    mem[5023] = 'd664;
    mem[5024] = 'd88;
    mem[5025] = 'd668;
    mem[5026] = 'd92;
    mem[5027] = 'd672;
    mem[5028] = 'd88;
    mem[5029] = 'd672;
    mem[5030] = 'd88;
    mem[5031] = 'd672;
    mem[5032] = 'd88;
    mem[5033] = 'd672;
    mem[5034] = 'd88;
    mem[5035] = 'd668;
    mem[5036] = 'd88;
    mem[5037] = 'd664;
    mem[5038] = 'd84;
    mem[5039] = 'd656;
    mem[5040] = 'd80;
    mem[5041] = 'd644;
    mem[5042] = 'd72;
    mem[5043] = 'd628;
    mem[5044] = 'd64;
    mem[5045] = 'd604;
    mem[5046] = 'd56;
    mem[5047] = 'd572;
    mem[5048] = 'd36;
    mem[5049] = 'd532;
    mem[5050] = 'd24;
    mem[5051] = 'd480;
    mem[5052] = 'd196;
    mem[5053] = 'd520;
    mem[5054] = 'd892;
    mem[5055] = 'd940;
    mem[5056] = 'd1012;
    mem[5057] = 'd1016;
    mem[5058] = 'd1016;
    mem[5059] = 'd1020;
    mem[5060] = 'd1020;
    mem[5061] = 'd1020;
    mem[5062] = 'd1020;
    mem[5063] = 'd1020;
    mem[5064] = 'd1020;
    mem[5065] = 'd1020;
    mem[5066] = 'd1020;
    mem[5067] = 'd1020;
    mem[5068] = 'd1020;
    mem[5069] = 'd1020;
    mem[5070] = 'd1020;
    mem[5071] = 'd1020;
    mem[5072] = 'd1020;
    mem[5073] = 'd1020;
    mem[5074] = 'd1020;
    mem[5075] = 'd1020;
    mem[5076] = 'd1020;
    mem[5077] = 'd1020;
    mem[5078] = 'd1020;
    mem[5079] = 'd1020;
    mem[5080] = 'd1020;
    mem[5081] = 'd1020;
    mem[5082] = 'd940;
    mem[5083] = 'd988;
    mem[5084] = 'd540;
    mem[5085] = 'd840;
    mem[5086] = 'd476;
    mem[5087] = 'd844;
    mem[5088] = 'd528;
    mem[5089] = 'd876;
    mem[5090] = 'd572;
    mem[5091] = 'd900;
    mem[5092] = 'd600;
    mem[5093] = 'd924;
    mem[5094] = 'd624;
    mem[5095] = 'd948;
    mem[5096] = 'd640;
    mem[5097] = 'd964;
    mem[5098] = 'd656;
    mem[5099] = 'd980;
    mem[5100] = 'd664;
    mem[5101] = 'd988;
    mem[5102] = 'd668;
    mem[5103] = 'd996;
    mem[5104] = 'd672;
    mem[5105] = 'd996;
    mem[5106] = 'd672;
    mem[5107] = 'd1000;
    mem[5108] = 'd672;
    mem[5109] = 'd1000;
    mem[5110] = 'd672;
    mem[5111] = 'd996;
    mem[5112] = 'd668;
    mem[5113] = 'd996;
    mem[5114] = 'd664;
    mem[5115] = 'd988;
    mem[5116] = 'd656;
    mem[5117] = 'd980;
    mem[5118] = 'd644;
    mem[5119] = 'd964;
    mem[5120] = 'd628;
    mem[5121] = 'd948;
    mem[5122] = 'd604;
    mem[5123] = 'd928;
    mem[5124] = 'd572;
    mem[5125] = 'd904;
    mem[5126] = 'd532;
    mem[5127] = 'd880;
    mem[5128] = 'd480;
    mem[5129] = 'd848;
    mem[5130] = 'd520;
    mem[5131] = 'd832;
    mem[5132] = 'd940;
    mem[5133] = 'd988;
    mem[5134] = 'd1016;
    mem[5135] = 'd1020;
    mem[5136] = 'd1020;
    mem[5137] = 'd1020;
    mem[5138] = 'd1020;
    mem[5139] = 'd1020;
    mem[5140] = 'd1020;
    mem[5141] = 'd1020;
    mem[5142] = 'd1020;
    mem[5143] = 'd1020;
    mem[5144] = 'd1020;
    mem[5145] = 'd1020;
    mem[5146] = 'd1020;
    mem[5147] = 'd1020;
    mem[5148] = 'd1020;
    mem[5149] = 'd1020;
    mem[5150] = 'd1020;
    mem[5151] = 'd1020;
    mem[5152] = 'd1020;
    mem[5153] = 'd1020;
    mem[5154] = 'd1020;
    mem[5155] = 'd1020;
    mem[5156] = 'd1020;
    mem[5157] = 'd1020;
    mem[5158] = 'd1016;
    mem[5159] = 'd1020;
    mem[5160] = 'd1012;
    mem[5161] = 'd1020;
    mem[5162] = 'd944;
    mem[5163] = 'd976;
    mem[5164] = 'd416;
    mem[5165] = 'd664;
    mem[5166] = 'd24;
    mem[5167] = 'd456;
    mem[5168] = 'd28;
    mem[5169] = 'd504;
    mem[5170] = 'd40;
    mem[5171] = 'd544;
    mem[5172] = 'd52;
    mem[5173] = 'd576;
    mem[5174] = 'd60;
    mem[5175] = 'd596;
    mem[5176] = 'd68;
    mem[5177] = 'd616;
    mem[5178] = 'd72;
    mem[5179] = 'd628;
    mem[5180] = 'd76;
    mem[5181] = 'd636;
    mem[5182] = 'd80;
    mem[5183] = 'd644;
    mem[5184] = 'd80;
    mem[5185] = 'd644;
    mem[5186] = 'd80;
    mem[5187] = 'd644;
    mem[5188] = 'd80;
    mem[5189] = 'd640;
    mem[5190] = 'd76;
    mem[5191] = 'd636;
    mem[5192] = 'd72;
    mem[5193] = 'd628;
    mem[5194] = 'd68;
    mem[5195] = 'd620;
    mem[5196] = 'd60;
    mem[5197] = 'd600;
    mem[5198] = 'd52;
    mem[5199] = 'd580;
    mem[5200] = 'd44;
    mem[5201] = 'd548;
    mem[5202] = 'd32;
    mem[5203] = 'd508;
    mem[5204] = 'd24;
    mem[5205] = 'd456;
    mem[5206] = 'd388;
    mem[5207] = 'd648;
    mem[5208] = 'd932;
    mem[5209] = 'd968;
    mem[5210] = 'd1012;
    mem[5211] = 'd1016;
    mem[5212] = 'd1016;
    mem[5213] = 'd1020;
    mem[5214] = 'd1020;
    mem[5215] = 'd1020;
    mem[5216] = 'd1020;
    mem[5217] = 'd1020;
    mem[5218] = 'd1020;
    mem[5219] = 'd1020;
    mem[5220] = 'd1020;
    mem[5221] = 'd1020;
    mem[5222] = 'd1020;
    mem[5223] = 'd1020;
    mem[5224] = 'd1020;
    mem[5225] = 'd1020;
    mem[5226] = 'd1020;
    mem[5227] = 'd1020;
    mem[5228] = 'd1020;
    mem[5229] = 'd1020;
    mem[5230] = 'd1020;
    mem[5231] = 'd1020;
    mem[5232] = 'd1020;
    mem[5233] = 'd1020;
    mem[5234] = 'd1020;
    mem[5235] = 'd1020;
    mem[5236] = 'd1020;
    mem[5237] = 'd1020;
    mem[5238] = 'd1020;
    mem[5239] = 'd1020;
    mem[5240] = 'd976;
    mem[5241] = 'd1000;
    mem[5242] = 'd664;
    mem[5243] = 'd888;
    mem[5244] = 'd456;
    mem[5245] = 'd824;
    mem[5246] = 'd504;
    mem[5247] = 'd864;
    mem[5248] = 'd544;
    mem[5249] = 'd888;
    mem[5250] = 'd576;
    mem[5251] = 'd908;
    mem[5252] = 'd596;
    mem[5253] = 'd924;
    mem[5254] = 'd616;
    mem[5255] = 'd944;
    mem[5256] = 'd628;
    mem[5257] = 'd952;
    mem[5258] = 'd636;
    mem[5259] = 'd964;
    mem[5260] = 'd644;
    mem[5261] = 'd964;
    mem[5262] = 'd644;
    mem[5263] = 'd968;
    mem[5264] = 'd644;
    mem[5265] = 'd968;
    mem[5266] = 'd640;
    mem[5267] = 'd968;
    mem[5268] = 'd636;
    mem[5269] = 'd964;
    mem[5270] = 'd628;
    mem[5271] = 'd956;
    mem[5272] = 'd620;
    mem[5273] = 'd944;
    mem[5274] = 'd600;
    mem[5275] = 'd928;
    mem[5276] = 'd580;
    mem[5277] = 'd912;
    mem[5278] = 'd548;
    mem[5279] = 'd892;
    mem[5280] = 'd508;
    mem[5281] = 'd868;
    mem[5282] = 'd456;
    mem[5283] = 'd828;
    mem[5284] = 'd648;
    mem[5285] = 'd884;
    mem[5286] = 'd968;
    mem[5287] = 'd1000;
    mem[5288] = 'd1016;
    mem[5289] = 'd1020;
    mem[5290] = 'd1020;
    mem[5291] = 'd1020;
    mem[5292] = 'd1020;
    mem[5293] = 'd1020;
    mem[5294] = 'd1020;
    mem[5295] = 'd1020;
    mem[5296] = 'd1020;
    mem[5297] = 'd1020;
    mem[5298] = 'd1020;
    mem[5299] = 'd1020;
    mem[5300] = 'd1020;
    mem[5301] = 'd1020;
    mem[5302] = 'd1020;
    mem[5303] = 'd1020;
    mem[5304] = 'd1020;
    mem[5305] = 'd1020;
    mem[5306] = 'd1020;
    mem[5307] = 'd1020;
    mem[5308] = 'd1020;
    mem[5309] = 'd1020;
    mem[5310] = 'd1020;
    mem[5311] = 'd1020;
    mem[5312] = 'd1020;
    mem[5313] = 'd1020;
    mem[5314] = 'd1020;
    mem[5315] = 'd1020;
    mem[5316] = 'd1016;
    mem[5317] = 'd1020;
    mem[5318] = 'd1012;
    mem[5319] = 'd1020;
    mem[5320] = 'd1004;
    mem[5321] = 'd1012;
    mem[5322] = 'd708;
    mem[5323] = 'd832;
    mem[5324] = 'd180;
    mem[5325] = 'd520;
    mem[5326] = 'd16;
    mem[5327] = 'd460;
    mem[5328] = 'd28;
    mem[5329] = 'd508;
    mem[5330] = 'd40;
    mem[5331] = 'd536;
    mem[5332] = 'd48;
    mem[5333] = 'd560;
    mem[5334] = 'd52;
    mem[5335] = 'd580;
    mem[5336] = 'd56;
    mem[5337] = 'd588;
    mem[5338] = 'd60;
    mem[5339] = 'd596;
    mem[5340] = 'd60;
    mem[5341] = 'd600;
    mem[5342] = 'd60;
    mem[5343] = 'd600;
    mem[5344] = 'd60;
    mem[5345] = 'd600;
    mem[5346] = 'd56;
    mem[5347] = 'd592;
    mem[5348] = 'd52;
    mem[5349] = 'd580;
    mem[5350] = 'd48;
    mem[5351] = 'd564;
    mem[5352] = 'd40;
    mem[5353] = 'd540;
    mem[5354] = 'd28;
    mem[5355] = 'd508;
    mem[5356] = 'd20;
    mem[5357] = 'd464;
    mem[5358] = 'd168;
    mem[5359] = 'd512;
    mem[5360] = 'd680;
    mem[5361] = 'd820;
    mem[5362] = 'd1000;
    mem[5363] = 'd1012;
    mem[5364] = 'd1012;
    mem[5365] = 'd1016;
    mem[5366] = 'd1016;
    mem[5367] = 'd1020;
    mem[5368] = 'd1020;
    mem[5369] = 'd1020;
    mem[5370] = 'd1020;
    mem[5371] = 'd1020;
    mem[5372] = 'd1020;
    mem[5373] = 'd1020;
    mem[5374] = 'd1020;
    mem[5375] = 'd1020;
    mem[5376] = 'd1020;
    mem[5377] = 'd1020;
    mem[5378] = 'd1020;
    mem[5379] = 'd1020;
    mem[5380] = 'd1020;
    mem[5381] = 'd1020;
    mem[5382] = 'd1020;
    mem[5383] = 'd1020;
    mem[5384] = 'd1020;
    mem[5385] = 'd1020;
    mem[5386] = 'd1020;
    mem[5387] = 'd1020;
    mem[5388] = 'd1020;
    mem[5389] = 'd1020;
    mem[5390] = 'd1020;
    mem[5391] = 'd1020;
    mem[5392] = 'd1020;
    mem[5393] = 'd1020;
    mem[5394] = 'd1020;
    mem[5395] = 'd1020;
    mem[5396] = 'd1020;
    mem[5397] = 'd1020;
    mem[5398] = 'd1012;
    mem[5399] = 'd1020;
    mem[5400] = 'd832;
    mem[5401] = 'd944;
    mem[5402] = 'd520;
    mem[5403] = 'd832;
    mem[5404] = 'd460;
    mem[5405] = 'd836;
    mem[5406] = 'd508;
    mem[5407] = 'd868;
    mem[5408] = 'd536;
    mem[5409] = 'd888;
    mem[5410] = 'd560;
    mem[5411] = 'd904;
    mem[5412] = 'd580;
    mem[5413] = 'd912;
    mem[5414] = 'd588;
    mem[5415] = 'd924;
    mem[5416] = 'd596;
    mem[5417] = 'd928;
    mem[5418] = 'd600;
    mem[5419] = 'd932;
    mem[5420] = 'd600;
    mem[5421] = 'd932;
    mem[5422] = 'd600;
    mem[5423] = 'd932;
    mem[5424] = 'd592;
    mem[5425] = 'd924;
    mem[5426] = 'd580;
    mem[5427] = 'd916;
    mem[5428] = 'd564;
    mem[5429] = 'd904;
    mem[5430] = 'd540;
    mem[5431] = 'd888;
    mem[5432] = 'd508;
    mem[5433] = 'd868;
    mem[5434] = 'd464;
    mem[5435] = 'd840;
    mem[5436] = 'd512;
    mem[5437] = 'd832;
    mem[5438] = 'd820;
    mem[5439] = 'd940;
    mem[5440] = 'd1012;
    mem[5441] = 'd1020;
    mem[5442] = 'd1016;
    mem[5443] = 'd1020;
    mem[5444] = 'd1020;
    mem[5445] = 'd1020;
    mem[5446] = 'd1020;
    mem[5447] = 'd1020;
    mem[5448] = 'd1020;
    mem[5449] = 'd1020;
    mem[5450] = 'd1020;
    mem[5451] = 'd1020;
    mem[5452] = 'd1020;
    mem[5453] = 'd1020;
    mem[5454] = 'd1020;
    mem[5455] = 'd1020;
    mem[5456] = 'd1020;
    mem[5457] = 'd1020;
    mem[5458] = 'd1020;
    mem[5459] = 'd1020;
    mem[5460] = 'd1020;
    mem[5461] = 'd1020;
    mem[5462] = 'd1020;
    mem[5463] = 'd1020;
    mem[5464] = 'd1020;
    mem[5465] = 'd1020;
    mem[5466] = 'd1020;
    mem[5467] = 'd1020;
    mem[5468] = 'd1020;
    mem[5469] = 'd1020;
    mem[5470] = 'd1020;
    mem[5471] = 'd1020;
    mem[5472] = 'd1020;
    mem[5473] = 'd1020;
    mem[5474] = 'd1020;
    mem[5475] = 'd1020;
    mem[5476] = 'd1016;
    mem[5477] = 'd1020;
    mem[5478] = 'd1008;
    mem[5479] = 'd1016;
    mem[5480] = 'd968;
    mem[5481] = 'd992;
    mem[5482] = 'd724;
    mem[5483] = 'd840;
    mem[5484] = 'd336;
    mem[5485] = 'd604;
    mem[5486] = 'd68;
    mem[5487] = 'd464;
    mem[5488] = 'd16;
    mem[5489] = 'd468;
    mem[5490] = 'd24;
    mem[5491] = 'd496;
    mem[5492] = 'd28;
    mem[5493] = 'd512;
    mem[5494] = 'd32;
    mem[5495] = 'd524;
    mem[5496] = 'd32;
    mem[5497] = 'd528;
    mem[5498] = 'd32;
    mem[5499] = 'd528;
    mem[5500] = 'd32;
    mem[5501] = 'd524;
    mem[5502] = 'd32;
    mem[5503] = 'd512;
    mem[5504] = 'd24;
    mem[5505] = 'd496;
    mem[5506] = 'd20;
    mem[5507] = 'd472;
    mem[5508] = 'd32;
    mem[5509] = 'd436;
    mem[5510] = 'd328;
    mem[5511] = 'd608;
    mem[5512] = 'd720;
    mem[5513] = 'd836;
    mem[5514] = 'd972;
    mem[5515] = 'd996;
    mem[5516] = 'd1008;
    mem[5517] = 'd1016;
    mem[5518] = 'd1012;
    mem[5519] = 'd1020;
    mem[5520] = 'd1016;
    mem[5521] = 'd1020;
    mem[5522] = 'd1020;
    mem[5523] = 'd1020;
    mem[5524] = 'd1020;
    mem[5525] = 'd1020;
    mem[5526] = 'd1020;
    mem[5527] = 'd1020;
    mem[5528] = 'd1020;
    mem[5529] = 'd1020;
    mem[5530] = 'd1020;
    mem[5531] = 'd1020;
    mem[5532] = 'd1020;
    mem[5533] = 'd1020;
    mem[5534] = 'd1020;
    mem[5535] = 'd1020;
    mem[5536] = 'd1020;
    mem[5537] = 'd1020;
    mem[5538] = 'd1020;
    mem[5539] = 'd1020;
    mem[5540] = 'd1020;
    mem[5541] = 'd1020;
    mem[5542] = 'd1020;
    mem[5543] = 'd1020;
    mem[5544] = 'd1020;
    mem[5545] = 'd1020;
    mem[5546] = 'd1020;
    mem[5547] = 'd1020;
    mem[5548] = 'd1020;
    mem[5549] = 'd1020;
    mem[5550] = 'd1020;
    mem[5551] = 'd1020;
    mem[5552] = 'd1020;
    mem[5553] = 'd1020;
    mem[5554] = 'd1020;
    mem[5555] = 'd1020;
    mem[5556] = 'd1016;
    mem[5557] = 'd1020;
    mem[5558] = 'd992;
    mem[5559] = 'd1008;
    mem[5560] = 'd840;
    mem[5561] = 'd952;
    mem[5562] = 'd604;
    mem[5563] = 'd856;
    mem[5564] = 'd464;
    mem[5565] = 'd816;
    mem[5566] = 'd468;
    mem[5567] = 'd840;
    mem[5568] = 'd496;
    mem[5569] = 'd860;
    mem[5570] = 'd512;
    mem[5571] = 'd872;
    mem[5572] = 'd524;
    mem[5573] = 'd876;
    mem[5574] = 'd528;
    mem[5575] = 'd880;
    mem[5576] = 'd528;
    mem[5577] = 'd880;
    mem[5578] = 'd524;
    mem[5579] = 'd876;
    mem[5580] = 'd512;
    mem[5581] = 'd872;
    mem[5582] = 'd496;
    mem[5583] = 'd860;
    mem[5584] = 'd472;
    mem[5585] = 'd840;
    mem[5586] = 'd436;
    mem[5587] = 'd804;
    mem[5588] = 'd608;
    mem[5589] = 'd860;
    mem[5590] = 'd836;
    mem[5591] = 'd948;
    mem[5592] = 'd996;
    mem[5593] = 'd1012;
    mem[5594] = 'd1016;
    mem[5595] = 'd1020;
    mem[5596] = 'd1020;
    mem[5597] = 'd1020;
    mem[5598] = 'd1020;
    mem[5599] = 'd1020;
    mem[5600] = 'd1020;
    mem[5601] = 'd1020;
    mem[5602] = 'd1020;
    mem[5603] = 'd1020;
    mem[5604] = 'd1020;
    mem[5605] = 'd1020;
    mem[5606] = 'd1020;
    mem[5607] = 'd1020;
    mem[5608] = 'd1020;
    mem[5609] = 'd1020;
    mem[5610] = 'd1020;
    mem[5611] = 'd1020;
    mem[5612] = 'd1020;
    mem[5613] = 'd1020;
    mem[5614] = 'd1020;
    mem[5615] = 'd1020;
    mem[5616] = 'd1020;
    mem[5617] = 'd1020;
    mem[5618] = 'd1020;
    mem[5619] = 'd1020;
    mem[5620] = 'd1020;
    mem[5621] = 'd1020;
    mem[5622] = 'd1020;
    mem[5623] = 'd1020;
    mem[5624] = 'd1020;
    mem[5625] = 'd1020;
    mem[5626] = 'd1020;
    mem[5627] = 'd1020;
    mem[5628] = 'd1020;
    mem[5629] = 'd1020;
    mem[5630] = 'd1020;
    mem[5631] = 'd1020;
    mem[5632] = 'd1020;
    mem[5633] = 'd1020;
    mem[5634] = 'd1016;
    mem[5635] = 'd1020;
    mem[5636] = 'd1012;
    mem[5637] = 'd1016;
    mem[5638] = 'd1012;
    mem[5639] = 'd1016;
    mem[5640] = 'd1008;
    mem[5641] = 'd1016;
    mem[5642] = 'd916;
    mem[5643] = 'd964;
    mem[5644] = 'd652;
    mem[5645] = 'd788;
    mem[5646] = 'd424;
    mem[5647] = 'd652;
    mem[5648] = 'd252;
    mem[5649] = 'd556;
    mem[5650] = 'd148;
    mem[5651] = 'd496;
    mem[5652] = 'd100;
    mem[5653] = 'd472;
    mem[5654] = 'd100;
    mem[5655] = 'd472;
    mem[5656] = 'd144;
    mem[5657] = 'd496;
    mem[5658] = 'd248;
    mem[5659] = 'd552;
    mem[5660] = 'd416;
    mem[5661] = 'd648;
    mem[5662] = 'd652;
    mem[5663] = 'd792;
    mem[5664] = 'd952;
    mem[5665] = 'd984;
    mem[5666] = 'd1004;
    mem[5667] = 'd1016;
    mem[5668] = 'd1012;
    mem[5669] = 'd1016;
    mem[5670] = 'd1016;
    mem[5671] = 'd1020;
    mem[5672] = 'd1016;
    mem[5673] = 'd1020;
    mem[5674] = 'd1020;
    mem[5675] = 'd1020;
    mem[5676] = 'd1020;
    mem[5677] = 'd1020;
    mem[5678] = 'd1020;
    mem[5679] = 'd1020;
    mem[5680] = 'd1020;
    mem[5681] = 'd1020;
    mem[5682] = 'd1020;
    mem[5683] = 'd1020;
    mem[5684] = 'd1020;
    mem[5685] = 'd1020;
    mem[5686] = 'd1020;
    mem[5687] = 'd1020;
    mem[5688] = 'd1020;
    mem[5689] = 'd1020;
    mem[5690] = 'd1020;
    mem[5691] = 'd1020;
    mem[5692] = 'd1020;
    mem[5693] = 'd1020;
    mem[5694] = 'd1020;
    mem[5695] = 'd1020;
    mem[5696] = 'd1020;
    mem[5697] = 'd1020;
    mem[5698] = 'd1020;
    mem[5699] = 'd1020;
    mem[5700] = 'd1020;
    mem[5701] = 'd1020;
    mem[5702] = 'd1020;
    mem[5703] = 'd1020;
    mem[5704] = 'd1020;
    mem[5705] = 'd1020;
    mem[5706] = 'd1020;
    mem[5707] = 'd1020;
    mem[5708] = 'd1020;
    mem[5709] = 'd1020;
    mem[5710] = 'd1020;
    mem[5711] = 'd1020;
    mem[5712] = 'd1020;
    mem[5713] = 'd1020;
    mem[5714] = 'd1016;
    mem[5715] = 'd1020;
    mem[5716] = 'd1016;
    mem[5717] = 'd1020;
    mem[5718] = 'd1016;
    mem[5719] = 'd1020;
    mem[5720] = 'd964;
    mem[5721] = 'd996;
    mem[5722] = 'd788;
    mem[5723] = 'd924;
    mem[5724] = 'd652;
    mem[5725] = 'd868;
    mem[5726] = 'd556;
    mem[5727] = 'd836;
    mem[5728] = 'd496;
    mem[5729] = 'd816;
    mem[5730] = 'd472;
    mem[5731] = 'd808;
    mem[5732] = 'd472;
    mem[5733] = 'd808;
    mem[5734] = 'd496;
    mem[5735] = 'd816;
    mem[5736] = 'd552;
    mem[5737] = 'd836;
    mem[5738] = 'd648;
    mem[5739] = 'd868;
    mem[5740] = 'd792;
    mem[5741] = 'd920;
    mem[5742] = 'd984;
    mem[5743] = 'd1008;
    mem[5744] = 'd1016;
    mem[5745] = 'd1020;
    mem[5746] = 'd1016;
    mem[5747] = 'd1020;
    mem[5748] = 'd1020;
    mem[5749] = 'd1020;
    mem[5750] = 'd1020;
    mem[5751] = 'd1020;
    mem[5752] = 'd1020;
    mem[5753] = 'd1020;
    mem[5754] = 'd1020;
    mem[5755] = 'd1020;
    mem[5756] = 'd1020;
    mem[5757] = 'd1020;
    mem[5758] = 'd1020;
    mem[5759] = 'd1020;
    mem[5760] = 'd1020;
    mem[5761] = 'd1020;
    mem[5762] = 'd1020;
    mem[5763] = 'd1020;
    mem[5764] = 'd1020;
    mem[5765] = 'd1020;
    mem[5766] = 'd1020;
    mem[5767] = 'd1020;
    mem[5768] = 'd1020;
    mem[5769] = 'd1020;
    mem[5770] = 'd1020;
    mem[5771] = 'd1020;
    mem[5772] = 'd1020;
    mem[5773] = 'd1020;
    mem[5774] = 'd1020;
    mem[5775] = 'd1020;
    mem[5776] = 'd1020;
    mem[5777] = 'd1020;
    mem[5778] = 'd1020;
    mem[5779] = 'd1020;
    mem[5780] = 'd1020;
    mem[5781] = 'd1020;
    mem[5782] = 'd1020;
    mem[5783] = 'd1020;
    mem[5784] = 'd1020;
    mem[5785] = 'd1020;
    mem[5786] = 'd1020;
    mem[5787] = 'd1020;
    mem[5788] = 'd1020;
    mem[5789] = 'd1020;
    mem[5790] = 'd1020;
    mem[5791] = 'd1020;
    mem[5792] = 'd1020;
    mem[5793] = 'd1020;
    mem[5794] = 'd1016;
    mem[5795] = 'd1020;
    mem[5796] = 'd1016;
    mem[5797] = 'd1020;
    mem[5798] = 'd1012;
    mem[5799] = 'd1016;
    mem[5800] = 'd1012;
    mem[5801] = 'd1016;
    mem[5802] = 'd1008;
    mem[5803] = 'd1016;
    mem[5804] = 'd1008;
    mem[5805] = 'd1016;
    mem[5806] = 'd1008;
    mem[5807] = 'd1016;
    mem[5808] = 'd1004;
    mem[5809] = 'd1012;
    mem[5810] = 'd1000;
    mem[5811] = 'd1012;
    mem[5812] = 'd1008;
    mem[5813] = 'd1016;
    mem[5814] = 'd1008;
    mem[5815] = 'd1016;
    mem[5816] = 'd1008;
    mem[5817] = 'd1016;
    mem[5818] = 'd1008;
    mem[5819] = 'd1016;
    mem[5820] = 'd1012;
    mem[5821] = 'd1016;
    mem[5822] = 'd1016;
    mem[5823] = 'd1020;
    mem[5824] = 'd1016;
    mem[5825] = 'd1020;
    mem[5826] = 'd1020;
    mem[5827] = 'd1020;
    mem[5828] = 'd1020;
    mem[5829] = 'd1020;
    mem[5830] = 'd1020;
    mem[5831] = 'd1020;
    mem[5832] = 'd1020;
    mem[5833] = 'd1020;
    mem[5834] = 'd1020;
    mem[5835] = 'd1020;
    mem[5836] = 'd1020;
    mem[5837] = 'd1020;
    mem[5838] = 'd1020;
    mem[5839] = 'd1020;
    mem[5840] = 'd1020;
    mem[5841] = 'd1020;
    mem[5842] = 'd1020;
    mem[5843] = 'd1020;
    mem[5844] = 'd1020;
    mem[5845] = 'd1020;
    mem[5846] = 'd1020;
    mem[5847] = 'd1020;
    mem[5848] = 'd1020;
    mem[5849] = 'd1020;
    mem[5850] = 'd1020;
    mem[5851] = 'd1020;
    mem[5852] = 'd1020;
    mem[5853] = 'd1020;
    mem[5854] = 'd1020;
    mem[5855] = 'd1020;
    mem[5856] = 'd1020;
    mem[5857] = 'd1020;
    mem[5858] = 'd1020;
    mem[5859] = 'd1020;
    mem[5860] = 'd1020;
    mem[5861] = 'd1020;
    mem[5862] = 'd1020;
    mem[5863] = 'd1020;
    mem[5864] = 'd1020;
    mem[5865] = 'd1020;
    mem[5866] = 'd1020;
    mem[5867] = 'd1020;
    mem[5868] = 'd1020;
    mem[5869] = 'd1020;
    mem[5870] = 'd1020;
    mem[5871] = 'd1020;
    mem[5872] = 'd1020;
    mem[5873] = 'd1020;
    mem[5874] = 'd1020;
    mem[5875] = 'd1020;
    mem[5876] = 'd1016;
    mem[5877] = 'd1020;
    mem[5878] = 'd1016;
    mem[5879] = 'd1020;
    mem[5880] = 'd1016;
    mem[5881] = 'd1020;
    mem[5882] = 'd1016;
    mem[5883] = 'd1020;
    mem[5884] = 'd1016;
    mem[5885] = 'd1020;
    mem[5886] = 'd1012;
    mem[5887] = 'd1020;
    mem[5888] = 'd1012;
    mem[5889] = 'd1020;
    mem[5890] = 'd1016;
    mem[5891] = 'd1020;
    mem[5892] = 'd1016;
    mem[5893] = 'd1020;
    mem[5894] = 'd1016;
    mem[5895] = 'd1020;
    mem[5896] = 'd1016;
    mem[5897] = 'd1020;
    mem[5898] = 'd1016;
    mem[5899] = 'd1020;
    mem[5900] = 'd1020;
    mem[5901] = 'd1020;
    mem[5902] = 'd1020;
    mem[5903] = 'd1020;
    mem[5904] = 'd1020;
    mem[5905] = 'd1020;
    mem[5906] = 'd1020;
    mem[5907] = 'd1020;
    mem[5908] = 'd1020;
    mem[5909] = 'd1020;
    mem[5910] = 'd1020;
    mem[5911] = 'd1020;
    mem[5912] = 'd1020;
    mem[5913] = 'd1020;
    mem[5914] = 'd1020;
    mem[5915] = 'd1020;
    mem[5916] = 'd1020;
    mem[5917] = 'd1020;
    mem[5918] = 'd1020;
    mem[5919] = 'd1020;
    mem[5920] = 'd1020;
    mem[5921] = 'd1020;
    mem[5922] = 'd1020;
    mem[5923] = 'd1020;
    mem[5924] = 'd1020;
    mem[5925] = 'd1020;
    mem[5926] = 'd1020;
    mem[5927] = 'd1020;

end

endmodule

module image_gen_colorbar #(
    parameter X_RESOLUTION = 1288,
    parameter Y_RESOLUTION = 768,
    parameter H_FRONT_PORCH = 50, // 2x X_RESOLUTION
    parameter H_BACK_PORCH = 50, // ~ 2.2x X_RESOLUTION
    parameter V_FRONT_PORCH = 2,
    parameter V_BACK_PORCH = 2,
    parameter H_SYNC_PULSE_WIDTH = 44,
    parameter V_SYNC_PULSE_WIDTH = 4
) (
    input logic pixel_clock_in,
    input logic reset_n_in,

    output logic [9:0] pixel_data_red_out,
    output logic [9:0] pixel_data_green_out,
    output logic [9:0] pixel_data_blue_out,
    output logic [9:0] pixel_data_out,

    output logic line_valid,
    output logic frame_valid
);

parameter H_START = H_SYNC_PULSE_WIDTH + H_BACK_PORCH;

logic [31:0] x_counter;
logic [31:0] y_counter;
logic [31:0] pixel_counter;

logic [9:0] mem[5927:0];

always @(posedge pixel_clock_in) begin

    if(!reset_n_in) begin

        pixel_data_red_out <= 0;
        pixel_data_green_out <= 0;
        pixel_data_blue_out <= 0;
        line_valid <= 0;
        frame_valid <= 0;

        x_counter <= 0;
        y_counter <= 0;
        pixel_counter <= 0;

    end 

    else begin
            
        // Increment counters
        if (x_counter <= (H_START + X_RESOLUTION + H_FRONT_PORCH)) begin
            x_counter <= x_counter + 1;
        end

        else begin
            x_counter <= 0;

            if (y_counter <= (V_SYNC_PULSE_WIDTH + V_BACK_PORCH + Y_RESOLUTION + V_FRONT_PORCH)) begin
                y_counter <= y_counter + 1;
            end

            else begin
                y_counter <= 0;
            end 

        end

        // Output line valud
        if ((x_counter >= (H_START)) &&
            (x_counter < (H_START + X_RESOLUTION)) &&
            (y_counter >= (V_SYNC_PULSE_WIDTH + V_BACK_PORCH)) &&
            (y_counter < (V_SYNC_PULSE_WIDTH + V_BACK_PORCH + Y_RESOLUTION))) begin
                
            line_valid <= 1;

            pixel_counter <= pixel_counter + 1;

            if ((x_counter >= (H_START)) &&
                (x_counter < (H_START + 100))) begin
                    pixel_data_red_out <= 'h3ff;
                    pixel_data_green_out <= 'h00;
                    pixel_data_blue_out <= 'h00;

                    if (!x_counter[0] && !y_counter[0]) pixel_data_out <= 'h0; //b
                    else if (x_counter[1] && !y_counter[0]) pixel_data_out <= 'h0; //g
                    else if (!x_counter[0] && y_counter[0]) pixel_data_out <= 'h0; //g
                    else if (x_counter[0] && y_counter[0]) pixel_data_out <= 'h3ff; //r
                end
            else if ((x_counter >= (H_START + 100)) &&
                (x_counter < (H_START + 200))) begin
                    pixel_data_red_out <= 'h00;
                    pixel_data_green_out <= 'h3ff;
                    pixel_data_blue_out <= 'h00;

                    if (!x_counter[0] && !y_counter[0]) pixel_data_out <= 'h3ff; //b
                    else if (x_counter[1] && !y_counter[0]) pixel_data_out <= 'h3ff; //g
                    else if (!x_counter[0] && y_counter[0]) pixel_data_out <= 'h3ff; //g
                    else if (x_counter[0] && y_counter[0]) pixel_data_out <= 'h0; //r
                end

            else if ((x_counter >= (H_START + 200)) &&
                (x_counter < (H_START + 300))) begin
                    pixel_data_red_out <= 'h00;
                    pixel_data_green_out <= 'h00;
                    pixel_data_blue_out <= 'h3ff;

                    if (!x_counter[0] && !y_counter[0]) pixel_data_out <= 'h3ff; //b
                    else if (x_counter[1] && !y_counter[0]) pixel_data_out <= 'h0; //g
                    else if (!x_counter[0] && y_counter[0]) pixel_data_out <= 'h0; //g
                    else if (x_counter[0] && y_counter[0]) pixel_data_out <= 'h0; //r
                end

            else if ((x_counter >= (H_START + 300)) &&
                (x_counter < (H_START + 400))) begin
                    pixel_data_red_out <= 'h3ff;
                    pixel_data_green_out <= 'h3ff;
                    pixel_data_blue_out <= 'h00;

                    if (!x_counter[0] && !y_counter[0]) pixel_data_out <= 'h0; //b
                    else if (x_counter[1] && !y_counter[0]) pixel_data_out <= 'h3ff; //g
                    else if (!x_counter[0] && y_counter[0]) pixel_data_out <= 'h3ff; //g
                    else if (x_counter[0] && y_counter[0]) pixel_data_out <= 'h3ff; //r
                end

            else if ((x_counter >= (H_START + 400)) &&
                (x_counter < (H_START + 500))) begin
                    pixel_data_red_out <= 'h00;
                    pixel_data_green_out <= 'h3ff;
                    pixel_data_blue_out <= 'h3ff;

                    if (!x_counter[0] && !y_counter[0]) pixel_data_out <= 'h0; //b
                    else if (x_counter[1] && !y_counter[0]) pixel_data_out <= 'h3ff; //g
                    else if (!x_counter[0] && y_counter[0]) pixel_data_out <= 'h3ff; //g
                    else if (x_counter[0] && y_counter[0]) pixel_data_out <= 'h0; //r
                end

            else if ((x_counter >= (H_START + 500)) &&
                (x_counter < (H_START + 600))) begin
                    pixel_data_red_out <= 'h3ff;
                    pixel_data_green_out <= 'h00;
                    pixel_data_blue_out <= 'h3ff;

                    if (!x_counter[0] && !y_counter[0]) pixel_data_out <= 'h3ff; //b
                    else if (x_counter[1] && !y_counter[0]) pixel_data_out <= 'h0; //g
                    else if (!x_counter[0] && y_counter[0]) pixel_data_out <= 'h0; //g
                    else if (x_counter[0] && y_counter[0]) pixel_data_out <= 'h3ff; //r
                end

            else begin
                    pixel_data_red_out <= 'h3ff;
                    pixel_data_green_out <= 'h3ff;
                    pixel_data_blue_out <= 'h3ff;

                    if (!x_counter[0] && !y_counter[0]) pixel_data_out <= 'h3ff; //b
                    else if (x_counter[1] && !y_counter[0]) pixel_data_out <= 'h3ff; //g
                    else if (!x_counter[0] && y_counter[0]) pixel_data_out <= 'h3ff; //g
                    else if (x_counter[0] && y_counter[0]) pixel_data_out <= 'h3ff; //r
                end

        end

        else begin
            line_valid <= 0;
        end

        // Output frame valid
        if (y_counter >= 0 &&
            y_counter < V_SYNC_PULSE_WIDTH) begin

            frame_valid <= 0;
            pixel_counter <= 0;

        end

        else begin
            frame_valid <= 1;
        end

    end

end

endmodule